module top(n0, n1, n2);
    input n0, n1;
    output n2;
    wire n0, n1;
    wire n2;
    wire [31:0] n3;
    wire [31:0] n4;
    wire [7:0] n5;
    wire n6, n7, n8, n9, n10, n11, n12, n13;
    wire n14, n15, n16, n17, n18, n19, n20, n21;
    wire n22, n23, n24, n25, n26, n27, n28, n29;
    wire n30, n31, n32, n33, n34, n35, n36, n37;
    wire n38, n39, n40, n41, n42, n43, n44, n45;
    wire n46, n47, n48, n49, n50, n51, n52, n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146, n147, n148, n149;
    wire n150, n151, n152, n153, n154, n155, n156, n157;
    wire n158, n159, n160, n161, n162, n163, n164, n165;
    wire n166, n167, n168, n169, n170, n171, n172, n173;
    wire n174, n175, n176, n177, n178, n179, n180, n181;
    wire n182, n183, n184, n185, n186, n187, n188, n189;
    wire n190, n191, n192, n193, n194, n195, n196, n197;
    wire n198, n199, n200, n201, n202, n203, n204, n205;
    wire n206, n207, n208, n209, n210, n211, n212, n213;
    wire n214, n215, n216, n217, n218, n219, n220, n221;
    wire n222, n223, n224, n225, n226, n227, n228, n229;
    wire n230, n231, n232, n233, n234, n235, n236, n237;
    wire n238, n239, n240, n241, n242, n243, n244, n245;
    wire n246, n247, n248, n249, n250, n251, n252, n253;
    wire n254, n255, n256, n257, n258, n259, n260, n261;
    wire n262, n263, n264, n265, n266, n267, n268, n269;
    wire n270, n271, n272, n273, n274, n275, n276, n277;
    wire n278, n279, n280, n281, n282, n283, n284, n285;
    wire n286, n287, n288, n289, n290, n291, n292, n293;
    wire n294, n295, n296, n297, n298, n299, n300, n301;
    wire n302, n303, n304, n305, n306, n307, n308, n309;
    wire n310, n311, n312, n313, n314, n315, n316, n317;
    wire n318, n319, n320, n321, n322, n323, n324, n325;
    wire n326, n327, n328, n329, n330, n331, n332, n333;
    wire n334, n335, n336, n337, n338, n339, n340, n341;
    wire n342, n343, n344, n345, n346, n347, n348, n349;
    wire n350, n351, n352, n353, n354, n355, n356, n357;
    wire n358, n359, n360, n361;
    not g0(n299 ,n335);
    dff g1(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n297), .Q(n3[1]));
    dff g2(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n298), .Q(n3[0]));
    dff g3(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n296), .Q(n3[2]));
    dff g4(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n295), .Q(n3[3]));
    or g5(n298 ,n279 ,n291);
    dff g6(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n290), .Q(n2));
    or g7(n297 ,n286 ,n294);
    or g8(n296 ,n285 ,n293);
    or g9(n295 ,n284 ,n292);
    dff g10(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n273), .Q(n4[1]));
    dff g11(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n282), .Q(n4[25]));
    dff g12(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n280), .Q(n4[26]));
    dff g13(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n288), .Q(n4[27]));
    dff g14(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n278), .Q(n4[28]));
    dff g15(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n277), .Q(n4[29]));
    dff g16(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n276), .Q(n4[30]));
    dff g17(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n268), .Q(n4[8]));
    dff g18(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n275), .Q(n4[31]));
    dff g19(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n283), .Q(n4[24]));
    dff g20(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n281), .Q(n4[23]));
    dff g21(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n272), .Q(n4[2]));
    dff g22(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n271), .Q(n4[3]));
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n287), .Q(n4[4]));
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n270), .Q(n4[5]));
    dff g25(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n269), .Q(n4[6]));
    dff g26(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n266), .Q(n4[7]));
    dff g27(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n251), .Q(n4[0]));
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n257), .Q(n4[18]));
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n265), .Q(n4[10]));
    dff g30(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n264), .Q(n4[11]));
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n263), .Q(n4[12]));
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n262), .Q(n4[13]));
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n261), .Q(n4[14]));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n260), .Q(n4[15]));
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n259), .Q(n4[16]));
    dff g36(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n258), .Q(n4[17]));
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n267), .Q(n4[9]));
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n256), .Q(n4[19]));
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n255), .Q(n4[20]));
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n254), .Q(n4[21]));
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n253), .Q(n4[22]));
    nor g42(n294 ,n215 ,n289);
    nor g43(n293 ,n218 ,n289);
    nor g44(n292 ,n207 ,n289);
    nor g45(n291 ,n3[0] ,n289);
    or g46(n290 ,n252 ,n274);
    nor g47(n288 ,n221 ,n247);
    nor g48(n287 ,n217 ,n247);
    nor g49(n286 ,n238 ,n248);
    nor g50(n285 ,n237 ,n248);
    nor g51(n284 ,n240 ,n248);
    nor g52(n283 ,n212 ,n247);
    nor g53(n282 ,n242 ,n247);
    nor g54(n281 ,n211 ,n247);
    nor g55(n280 ,n210 ,n247);
    nor g56(n279 ,n236 ,n248);
    nor g57(n278 ,n220 ,n247);
    nor g58(n277 ,n222 ,n247);
    nor g59(n276 ,n205 ,n247);
    nor g60(n275 ,n204 ,n247);
    nor g61(n274 ,n202 ,n247);
    nor g62(n273 ,n209 ,n247);
    nor g63(n272 ,n219 ,n247);
    nor g64(n271 ,n213 ,n247);
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n249), .Q(n337));
    or g66(n289 ,n299 ,n250);
    nor g67(n270 ,n225 ,n247);
    nor g68(n269 ,n208 ,n247);
    nor g69(n268 ,n203 ,n247);
    nor g70(n267 ,n235 ,n247);
    nor g71(n266 ,n206 ,n247);
    nor g72(n265 ,n229 ,n247);
    nor g73(n264 ,n234 ,n247);
    nor g74(n263 ,n223 ,n247);
    nor g75(n262 ,n216 ,n247);
    nor g76(n261 ,n227 ,n247);
    nor g77(n260 ,n214 ,n247);
    nor g78(n259 ,n226 ,n247);
    nor g79(n258 ,n231 ,n247);
    nor g80(n257 ,n224 ,n247);
    nor g81(n256 ,n233 ,n247);
    nor g82(n255 ,n228 ,n247);
    nor g83(n254 ,n232 ,n247);
    nor g84(n253 ,n230 ,n247);
    nor g85(n252 ,n241 ,n246);
    nor g86(n251 ,n4[0] ,n247);
    or g87(n250 ,n239 ,n245);
    nor g88(n249 ,n244 ,n245);
    not g89(n247 ,n246);
    or g90(n248 ,n337 ,n245);
    nor g91(n246 ,n243 ,n245);
    or g92(n245 ,n1 ,n6);
    not g93(n244 ,n243);
    nor g94(n243 ,n336 ,n327);
    not g95(n242 ,n324);
    not g96(n241 ,n2);
    not g97(n240 ,n3[3]);
    not g98(n239 ,n337);
    not g99(n238 ,n3[1]);
    not g100(n237 ,n3[2]);
    not g101(n236 ,n3[0]);
    not g102(n235 ,n308);
    not g103(n234 ,n310);
    not g104(n233 ,n318);
    not g105(n232 ,n320);
    not g106(n231 ,n316);
    not g107(n230 ,n321);
    not g108(n229 ,n309);
    not g109(n228 ,n319);
    not g110(n227 ,n313);
    not g111(n226 ,n315);
    not g112(n225 ,n304);
    not g113(n224 ,n317);
    not g114(n223 ,n311);
    not g115(n222 ,n331);
    not g116(n221 ,n329);
    not g117(n220 ,n330);
    not g118(n219 ,n301);
    not g119(n218 ,n333);
    not g120(n217 ,n303);
    not g121(n216 ,n312);
    not g122(n215 ,n332);
    not g123(n214 ,n314);
    not g124(n213 ,n302);
    not g125(n212 ,n323);
    not g126(n211 ,n322);
    not g127(n210 ,n328);
    not g128(n209 ,n300);
    not g129(n208 ,n305);
    not g130(n207 ,n334);
    not g131(n206 ,n306);
    not g132(n205 ,n325);
    not g133(n204 ,n326);
    not g134(n203 ,n307);
    not g135(n202 ,n336);
    xor g136(n326 ,n4[31] ,n114);
    nor g137(n325 ,n113 ,n114);
    nor g138(n114 ,n37 ,n112);
    nor g139(n113 ,n4[30] ,n111);
    xor g140(n331 ,n4[29] ,n109);
    not g141(n112 ,n111);
    nor g142(n111 ,n24 ,n110);
    nor g143(n330 ,n108 ,n109);
    not g144(n110 ,n109);
    nor g145(n109 ,n35 ,n107);
    nor g146(n108 ,n4[28] ,n106);
    xor g147(n329 ,n4[27] ,n104);
    not g148(n107 ,n106);
    nor g149(n106 ,n10 ,n105);
    nor g150(n328 ,n103 ,n104);
    xor g151(n324 ,n4[25] ,n102);
    not g152(n105 ,n104);
    nor g153(n104 ,n22 ,n101);
    nor g154(n103 ,n4[26] ,n100);
    nor g155(n323 ,n99 ,n102);
    nor g156(n102 ,n20 ,n98);
    not g157(n101 ,n100);
    nor g158(n100 ,n43 ,n98);
    nor g159(n99 ,n4[24] ,n97);
    xor g160(n322 ,n4[23] ,n95);
    not g161(n98 ,n97);
    nor g162(n97 ,n9 ,n96);
    nor g163(n321 ,n94 ,n95);
    xor g164(n320 ,n4[21] ,n93);
    xor g165(n318 ,n4[19] ,n92);
    not g166(n96 ,n95);
    nor g167(n95 ,n36 ,n91);
    nor g168(n94 ,n4[22] ,n90);
    nor g169(n319 ,n89 ,n93);
    nor g170(n317 ,n88 ,n92);
    xor g171(n316 ,n4[17] ,n87);
    nor g172(n93 ,n31 ,n84);
    nor g173(n92 ,n19 ,n86);
    not g174(n91 ,n90);
    nor g175(n90 ,n46 ,n84);
    nor g176(n89 ,n4[20] ,n83);
    nor g177(n88 ,n4[18] ,n85);
    nor g178(n315 ,n82 ,n87);
    nor g179(n87 ,n15 ,n81);
    not g180(n86 ,n85);
    nor g181(n85 ,n44 ,n81);
    not g182(n84 ,n83);
    nor g183(n83 ,n54 ,n81);
    nor g184(n82 ,n4[16] ,n80);
    xor g185(n314 ,n4[15] ,n78);
    not g186(n81 ,n80);
    nor g187(n80 ,n30 ,n79);
    nor g188(n313 ,n77 ,n78);
    xor g189(n312 ,n4[13] ,n76);
    xor g190(n310 ,n4[11] ,n75);
    or g191(n79 ,n13 ,n74);
    nor g192(n78 ,n30 ,n74);
    nor g193(n77 ,n4[14] ,n73);
    nor g194(n311 ,n71 ,n76);
    nor g195(n309 ,n72 ,n75);
    xor g196(n308 ,n4[9] ,n70);
    nor g197(n76 ,n18 ,n69);
    nor g198(n75 ,n16 ,n67);
    not g199(n74 ,n73);
    nor g200(n73 ,n45 ,n69);
    nor g201(n72 ,n4[10] ,n66);
    nor g202(n71 ,n4[12] ,n68);
    nor g203(n307 ,n65 ,n70);
    nor g204(n70 ,n25 ,n64);
    not g205(n69 ,n68);
    nor g206(n68 ,n55 ,n64);
    not g207(n67 ,n66);
    nor g208(n66 ,n42 ,n64);
    nor g209(n65 ,n4[8] ,n63);
    xor g210(n306 ,n4[7] ,n62);
    not g211(n64 ,n63);
    nor g212(n63 ,n27 ,n61);
    nor g213(n305 ,n60 ,n62);
    xor g214(n304 ,n4[5] ,n59);
    nor g215(n62 ,n27 ,n58);
    or g216(n61 ,n23 ,n58);
    nor g217(n60 ,n4[6] ,n57);
    nor g218(n303 ,n56 ,n59);
    nor g219(n59 ,n12 ,n53);
    not g220(n58 ,n57);
    nor g221(n57 ,n41 ,n53);
    nor g222(n56 ,n4[4] ,n52);
    xor g223(n302 ,n4[3] ,n50);
    or g224(n55 ,n16 ,n48);
    or g225(n54 ,n19 ,n51);
    not g226(n53 ,n52);
    nor g227(n52 ,n7 ,n49);
    nor g228(n301 ,n47 ,n50);
    or g229(n51 ,n14 ,n44);
    nor g230(n50 ,n32 ,n40);
    or g231(n49 ,n32 ,n40);
    or g232(n48 ,n11 ,n42);
    nor g233(n47 ,n4[2] ,n39);
    nor g234(n300 ,n39 ,n38);
    or g235(n46 ,n26 ,n31);
    or g236(n45 ,n8 ,n18);
    or g237(n44 ,n33 ,n15);
    or g238(n43 ,n17 ,n20);
    or g239(n42 ,n28 ,n25);
    or g240(n41 ,n29 ,n12);
    not g241(n40 ,n39);
    nor g242(n39 ,n21 ,n34);
    nor g243(n38 ,n4[1] ,n4[0]);
    not g244(n37 ,n4[30]);
    not g245(n36 ,n4[22]);
    not g246(n35 ,n4[28]);
    not g247(n34 ,n4[0]);
    not g248(n33 ,n4[17]);
    not g249(n32 ,n4[2]);
    not g250(n31 ,n4[20]);
    not g251(n30 ,n4[14]);
    not g252(n29 ,n4[5]);
    not g253(n28 ,n4[9]);
    not g254(n27 ,n4[6]);
    not g255(n26 ,n4[21]);
    not g256(n25 ,n4[8]);
    not g257(n24 ,n4[29]);
    not g258(n23 ,n4[7]);
    not g259(n22 ,n4[26]);
    not g260(n21 ,n4[1]);
    not g261(n20 ,n4[24]);
    not g262(n19 ,n4[18]);
    not g263(n18 ,n4[12]);
    not g264(n17 ,n4[25]);
    not g265(n16 ,n4[10]);
    not g266(n15 ,n4[16]);
    not g267(n14 ,n4[19]);
    not g268(n13 ,n4[15]);
    not g269(n12 ,n4[4]);
    not g270(n11 ,n4[11]);
    not g271(n10 ,n4[27]);
    not g272(n9 ,n4[23]);
    not g273(n8 ,n4[13]);
    not g274(n7 ,n4[3]);
    xor g275(n334 ,n3[3] ,n122);
    nor g276(n333 ,n121 ,n122);
    nor g277(n122 ,n117 ,n120);
    nor g278(n121 ,n3[2] ,n119);
    nor g279(n332 ,n119 ,n118);
    not g280(n120 ,n119);
    nor g281(n119 ,n115 ,n116);
    nor g282(n118 ,n3[1] ,n3[0]);
    not g283(n117 ,n3[2]);
    not g284(n116 ,n3[0]);
    not g285(n115 ,n3[1]);
    nor g286(n152 ,n148 ,n151);
    or g287(n151 ,n150 ,n149);
    or g288(n150 ,n137 ,n145);
    or g289(n149 ,n147 ,n146);
    or g290(n148 ,n142 ,n140);
    or g291(n147 ,n143 ,n141);
    or g292(n146 ,n139 ,n138);
    or g293(n145 ,n4[4] ,n144);
    nor g294(n144 ,n123 ,n130);
    or g295(n143 ,n136 ,n134);
    or g296(n142 ,n129 ,n135);
    or g297(n141 ,n132 ,n124);
    or g298(n140 ,n127 ,n131);
    or g299(n139 ,n128 ,n133);
    or g300(n138 ,n126 ,n125);
    or g301(n137 ,n4[6] ,n4[5]);
    or g302(n136 ,n4[30] ,n4[29]);
    or g303(n135 ,n4[12] ,n4[11]);
    or g304(n134 ,n4[28] ,n4[27]);
    or g305(n133 ,n4[20] ,n4[19]);
    or g306(n132 ,n4[26] ,n4[25]);
    or g307(n131 ,n4[8] ,n4[7]);
    nor g308(n130 ,n4[2] ,n4[1]);
    or g309(n129 ,n4[14] ,n4[13]);
    or g310(n128 ,n4[22] ,n4[21]);
    or g311(n127 ,n4[10] ,n4[9]);
    or g312(n126 ,n4[18] ,n4[17]);
    or g313(n125 ,n4[16] ,n4[15]);
    or g314(n124 ,n4[24] ,n4[23]);
    not g315(n123 ,n4[3]);
    or g316(n335 ,n153 ,n154);
    nor g317(n154 ,n3[2] ,n3[1]);
    not g318(n153 ,n3[3]);
    or g319(n336 ,n4[31] ,n201);
    nor g320(n201 ,n197 ,n200);
    or g321(n200 ,n190 ,n199);
    or g322(n199 ,n193 ,n198);
    or g323(n198 ,n181 ,n196);
    nor g324(n197 ,n180 ,n194);
    or g325(n196 ,n174 ,n195);
    or g326(n195 ,n173 ,n192);
    nor g327(n194 ,n176 ,n191);
    or g328(n193 ,n168 ,n187);
    or g329(n192 ,n4[25] ,n189);
    or g330(n191 ,n175 ,n188);
    or g331(n190 ,n182 ,n185);
    or g332(n189 ,n4[24] ,n184);
    nor g333(n188 ,n3[0] ,n186);
    or g334(n187 ,n4[4] ,n183);
    or g335(n186 ,n161 ,n178);
    or g336(n185 ,n172 ,n179);
    or g337(n184 ,n162 ,n169);
    or g338(n183 ,n167 ,n166);
    or g339(n182 ,n165 ,n163);
    or g340(n181 ,n164 ,n170);
    or g341(n180 ,n177 ,n171);
    or g342(n179 ,n4[12] ,n4[11]);
    nor g343(n178 ,n159 ,n4[1]);
    nor g344(n177 ,n160 ,n4[3]);
    nor g345(n176 ,n158 ,n3[2]);
    nor g346(n175 ,n156 ,n3[1]);
    nor g347(n174 ,n155 ,n3[3]);
    or g348(n173 ,n4[26] ,n4[23]);
    or g349(n172 ,n4[14] ,n4[13]);
    nor g350(n171 ,n157 ,n4[2]);
    or g351(n170 ,n4[28] ,n4[27]);
    or g352(n169 ,n4[20] ,n4[19]);
    or g353(n168 ,n4[6] ,n4[5]);
    or g354(n167 ,n4[10] ,n4[9]);
    or g355(n166 ,n4[8] ,n4[7]);
    or g356(n165 ,n4[18] ,n4[17]);
    or g357(n164 ,n4[30] ,n4[29]);
    or g358(n163 ,n4[16] ,n4[15]);
    or g359(n162 ,n4[22] ,n4[21]);
    not g360(n161 ,n4[0]);
    not g361(n160 ,n3[3]);
    not g362(n159 ,n3[1]);
    not g363(n158 ,n4[2]);
    not g364(n157 ,n3[2]);
    not g365(n156 ,n4[1]);
    not g366(n155 ,n4[3]);
    buf g367(n327 ,n152);
    dff g368(.RN(n338), .SN(1'b1), .CK(n0), .D(n361), .Q(n6));
    nor g369(n361 ,n360 ,n359);
    or g370(n360 ,n355 ,n358);
    or g371(n359 ,n356 ,n357);
    or g372(n358 ,n353 ,n352);
    or g373(n357 ,n354 ,n349);
    or g374(n356 ,n348 ,n347);
    or g375(n355 ,n351 ,n350);
    dff g376(.RN(n338), .SN(1'b1), .CK(n0), .D(n4[4]), .Q(n5[4]));
    dff g377(.RN(n338), .SN(1'b1), .CK(n0), .D(n4[1]), .Q(n5[1]));
    dff g378(.RN(n338), .SN(1'b1), .CK(n0), .D(n4[2]), .Q(n5[2]));
    dff g379(.RN(n338), .SN(1'b1), .CK(n0), .D(n4[3]), .Q(n5[3]));
    dff g380(.RN(n338), .SN(1'b1), .CK(n0), .D(n4[0]), .Q(n5[0]));
    dff g381(.RN(n338), .SN(1'b1), .CK(n0), .D(n4[5]), .Q(n5[5]));
    dff g382(.RN(n338), .SN(1'b1), .CK(n0), .D(n4[7]), .Q(n5[7]));
    dff g383(.RN(n338), .SN(1'b1), .CK(n0), .D(n4[6]), .Q(n5[6]));
    or g384(n354 ,n4[5] ,n4[3]);
    or g385(n353 ,n342 ,n341);
    or g386(n352 ,n339 ,n340);
    or g387(n351 ,n343 ,n346);
    or g388(n350 ,n345 ,n344);
    or g389(n349 ,n4[7] ,n4[1]);
    or g390(n348 ,n5[0] ,n5[2]);
    or g391(n347 ,n5[4] ,n5[6]);
    not g392(n346 ,n5[3]);
    not g393(n345 ,n5[5]);
    not g394(n344 ,n5[7]);
    not g395(n343 ,n5[1]);
    not g396(n342 ,n4[6]);
    not g397(n341 ,n4[4]);
    not g398(n340 ,n4[0]);
    not g399(n339 ,n4[2]);
    not g400(n338 ,n1);
endmodule
