module top(n0, n1, n2, n3);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3;
    wire [7:0] n4;
    wire [7:0] n5;
    wire [63:0] n6;
    wire [7:0] n7;
    wire [3:0] n8;
    wire [3:0] n9;
    wire [15:0] n10;
    wire [7:0] n11;
    wire [3:0] n12;
    wire [15:0] n13;
    wire [31:0] n14;
    wire [15:0] n15;
    wire [63:0] n16;
    wire [19:0] n17;
    wire n18, n19, n20, n21, n22, n23, n24, n25;
    wire n26, n27, n28, n29, n30, n31, n32, n33;
    wire n34, n35, n36, n37, n38, n39, n40, n41;
    wire n42, n43, n44, n45, n46, n47, n48, n49;
    wire n50, n51, n52, n53, n54, n55, n56, n57;
    wire n58, n59, n60, n61, n62, n63, n64, n65;
    wire n66, n67, n68, n69, n70, n71, n72, n73;
    wire n74, n75, n76, n77, n78, n79, n80, n81;
    wire n82, n83, n84, n85, n86, n87, n88, n89;
    wire n90, n91, n92, n93, n94, n95, n96, n97;
    wire n98, n99, n100, n101, n102, n103, n104, n105;
    wire n106, n107, n108, n109, n110, n111, n112, n113;
    wire n114, n115, n116, n117, n118, n119, n120, n121;
    wire n122, n123, n124, n125, n126, n127, n128, n129;
    wire n130, n131, n132, n133, n134, n135, n136, n137;
    wire n138, n139, n140, n141, n142, n143, n144, n145;
    wire n146, n147, n148, n149, n150, n151, n152, n153;
    wire n154, n155, n156, n157, n158, n159, n160, n161;
    wire n162, n163, n164, n165, n166, n167, n168, n169;
    wire n170, n171, n172, n173, n174, n175, n176, n177;
    wire n178, n179, n180, n181, n182, n183, n184, n185;
    wire n186, n187, n188, n189, n190, n191, n192, n193;
    wire n194, n195, n196, n197, n198, n199, n200, n201;
    wire n202, n203, n204, n205, n206, n207, n208, n209;
    wire n210, n211, n212, n213, n214, n215, n216, n217;
    wire n218, n219, n220, n221, n222, n223, n224, n225;
    wire n226, n227, n228, n229, n230, n231, n232, n233;
    wire n234, n235, n236, n237, n238, n239, n240, n241;
    wire n242, n243, n244, n245, n246, n247, n248, n249;
    wire n250, n251, n252, n253, n254, n255, n256, n257;
    wire n258, n259, n260, n261, n262, n263, n264, n265;
    wire n266, n267, n268, n269, n270, n271, n272, n273;
    wire n274, n275, n276, n277, n278, n279, n280, n281;
    wire n282, n283, n284, n285, n286, n287, n288, n289;
    wire n290, n291, n292, n293, n294, n295, n296, n297;
    wire n298, n299, n300, n301, n302, n303, n304, n305;
    wire n306, n307, n308, n309, n310, n311, n312, n313;
    wire n314, n315, n316, n317, n318, n319, n320, n321;
    wire n322, n323, n324, n325, n326, n327, n328, n329;
    wire n330, n331, n332, n333, n334, n335, n336, n337;
    wire n338, n339, n340, n341, n342, n343, n344, n345;
    wire n346, n347, n348, n349, n350, n351, n352, n353;
    wire n354, n355, n356, n357, n358, n359, n360, n361;
    wire n362, n363, n364, n365, n366, n367, n368, n369;
    wire n370, n371, n372, n373, n374, n375, n376, n377;
    wire n378, n379, n380, n381, n382, n383, n384, n385;
    wire n386, n387, n388, n389, n390, n391, n392, n393;
    wire n394, n395, n396, n397, n398, n399, n400, n401;
    wire n402, n403, n404, n405, n406, n407, n408, n409;
    wire n410, n411, n412, n413, n414, n415, n416, n417;
    wire n418, n419, n420, n421, n422, n423, n424, n425;
    wire n426, n427, n428, n429, n430, n431, n432, n433;
    wire n434, n435, n436, n437, n438, n439, n440, n441;
    wire n442, n443, n444, n445, n446, n447, n448, n449;
    wire n450, n451, n452, n453, n454, n455, n456, n457;
    wire n458, n459, n460, n461, n462, n463, n464, n465;
    wire n466, n467, n468, n469, n470, n471, n472, n473;
    wire n474, n475, n476, n477, n478, n479, n480, n481;
    wire n482, n483, n484, n485, n486, n487, n488, n489;
    wire n490, n491, n492, n493, n494, n495, n496, n497;
    wire n498, n499, n500, n501, n502, n503, n504, n505;
    wire n506, n507, n508, n509, n510, n511, n512, n513;
    wire n514, n515, n516, n517, n518, n519, n520, n521;
    wire n522, n523, n524, n525, n526, n527, n528, n529;
    wire n530, n531, n532, n533, n534, n535, n536, n537;
    wire n538, n539, n540, n541, n542, n543, n544, n545;
    wire n546, n547, n548, n549, n550, n551, n552, n553;
    wire n554, n555, n556, n557, n558, n559, n560, n561;
    wire n562, n563, n564, n565, n566, n567, n568, n569;
    wire n570, n571, n572, n573, n574, n575, n576, n577;
    nor g0(n302 ,n11[0] ,n11[1]);
    nor g1(n101 ,n78 ,n99);
    dff g2(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n387), .Q(n15[15]));
    or g3(n23 ,n15[4] ,n15[3]);
    or g4(n328 ,n246 ,n252);
    dff g5(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n572), .Q(n16[7]));
    not g6(n538 ,n17[15]);
    xnor g7(n333 ,n9[0] ,n16[7]);
    nor g8(n565 ,n538 ,n1);
    nor g9(n360 ,n321 ,n287);
    or g10(n48 ,n41 ,n42);
    nor g11(n344 ,n318 ,n298);
    not g12(n117 ,n116);
    dff g13(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n467), .Q(n11[2]));
    buf g14(n3[30], n3[31]);
    not g15(n158 ,n157);
    buf g16(n3[61], n3[63]);
    not g17(n239 ,n519);
    dff g18(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n477), .Q(n6[24]));
    nor g19(n296 ,n241 ,n498);
    xor g20(n572 ,n17[0] ,n2[0]);
    nor g21(n112 ,n15[9] ,n110);
    nor g22(n32 ,n20 ,n31);
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n281), .Q(n14[0]));
    xnor g24(n3[7] ,n491 ,n6[0]);
    nor g25(n466 ,n203 ,n453);
    nor g26(n306 ,n250 ,n193);
    dff g27(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n365), .Q(n10[9]));
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n363), .Q(n10[2]));
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n346), .Q(n10[15]));
    nor g30(n162 ,n10[7] ,n160);
    not g31(n134 ,n10[5]);
    or g32(n41 ,n10[13] ,n10[12]);
    or g33(n553 ,n17[5] ,n1);
    not g34(n39 ,n10[7]);
    nor g35(n301 ,n193 ,n11[0]);
    not g36(n497 ,n520);
    or g37(n472 ,n445 ,n462);
    or g38(n26 ,n15[11] ,n15[10]);
    not g39(n204 ,n16[55]);
    nor g40(n157 ,n134 ,n155);
    nor g41(n377 ,n233 ,n332);
    or g42(n332 ,n193 ,n197);
    nor g43(n562 ,n539 ,n1);
    buf g44(n3[5], n3[7]);
    nor g45(n465 ,n201 ,n453);
    nor g46(n191 ,n12[2] ,n189);
    not g47(n262 ,n15[8]);
    nor g48(n174 ,n10[11] ,n172);
    or g49(n419 ,n242 ,n380);
    nor g50(n323 ,n261 ,n194);
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n401), .Q(n15[0]));
    not g52(n259 ,n15[9]);
    not g53(n243 ,n11[2]);
    nor g54(n528 ,n112 ,n113);
    not g55(n186 ,n12[0]);
    nor g56(n501 ,n145 ,n144);
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n554), .Q(n17[15]));
    not g58(n120 ,n119);
    not g59(n544 ,n17[10]);
    nor g60(n294 ,n218 ,n498);
    not g61(n251 ,n12[3]);
    or g62(n554 ,n17[16] ,n1);
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n305), .Q(n5[4]));
    not g64(n90 ,n89);
    nor g65(n384 ,n193 ,n337);
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n405), .Q(n8[1]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n379), .Q(n10[14]));
    nor g68(n115 ,n15[10] ,n113);
    nor g69(n107 ,n80 ,n105);
    not g70(n161 ,n160);
    not g71(n218 ,n528);
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n394), .Q(n15[8]));
    buf g73(n3[41], n3[47]);
    not g74(n40 ,n10[6]);
    nor g75(n70 ,n64 ,n68);
    nor g76(n351 ,n323 ,n289);
    nor g77(n413 ,n240 ,n361);
    or g78(n380 ,n278 ,n357);
    nor g79(n424 ,n381 ,n411);
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n431), .Q(n12[3]));
    xnor g81(n481 ,n11[0] ,n12[0]);
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n471), .Q(n6[48]));
    not g83(n200 ,n16[39]);
    nor g84(n28 ,n19 ,n21);
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n366), .Q(n10[5]));
    nor g86(n518 ,n191 ,n192);
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n476), .Q(n6[16]));
    nor g88(n144 ,n10[1] ,n10[0]);
    nor g89(n510 ,n171 ,n172);
    buf g90(n3[8], n3[15]);
    nor g91(n324 ,n258 ,n194);
    or g92(n484 ,n4[0] ,n500);
    or g93(n477 ,n447 ,n466);
    or g94(n359 ,n196 ,n273);
    buf g95(n3[21], n3[23]);
    or g96(n60 ,n15[13] ,n15[12]);
    buf g97(n3[20], n3[23]);
    not g98(n114 ,n113);
    not g99(n255 ,n15[7]);
    xnor g100(n3[15] ,n491 ,n6[8]);
    nor g101(n369 ,n497 ,n300);
    nor g102(n416 ,n408 ,n414);
    not g103(n267 ,n5[5]);
    buf g104(n3[62], n3[63]);
    nor g105(n405 ,n193 ,n339);
    or g106(n470 ,n443 ,n460);
    xnor g107(n567 ,n17[7] ,n17[0]);
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n386), .Q(n9[0]));
    nor g109(n314 ,n255 ,n194);
    nor g110(n372 ,n215 ,n332);
    buf g111(n3[53], n3[55]);
    nor g112(n110 ,n79 ,n108);
    nor g113(n336 ,n311 ,n291);
    buf g114(n3[49], n3[55]);
    nor g115(n462 ,n206 ,n453);
    not g116(n257 ,n5[6]);
    not g117(n492 ,n5[3]);
    not g118(n146 ,n145);
    not g119(n135 ,n10[8]);
    nor g120(n448 ,n16[7] ,n441);
    not g121(n246 ,n12[0]);
    not g122(n201 ,n16[23]);
    nor g123(n435 ,n330 ,n419);
    not g124(n57 ,n15[5]);
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n389), .Q(n15[13]));
    buf g126(n3[0], n3[7]);
    not g127(n237 ,n535);
    nor g128(n119 ,n83 ,n117);
    not g129(n203 ,n16[31]);
    not g130(n248 ,n10[0]);
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n425), .Q(n8[2]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n552), .Q(n17[16]));
    nor g133(n156 ,n10[5] ,n154);
    xor g134(n517 ,n12[3] ,n192);
    or g135(n453 ,n193 ,n440);
    nor g136(n365 ,n227 ,n332);
    nor g137(n309 ,n193 ,n197);
    nor g138(n388 ,n193 ,n342);
    nor g139(n564 ,n546 ,n1);
    nor g140(n366 ,n208 ,n332);
    nor g141(n357 ,n244 ,n326);
    not g142(n252 ,n12[1]);
    not g143(n86 ,n15[0]);
    nor g144(n184 ,n140 ,n182);
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n307), .Q(n4[2]));
    not g146(n236 ,n2[2]);
    not g147(n108 ,n107);
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n561), .Q(n17[10]));
    not g149(n35 ,n10[5]);
    nor g150(n350 ,n327 ,n272);
    not g151(n87 ,n15[12]);
    or g152(n65 ,n15[3] ,n63);
    or g153(n72 ,n15[14] ,n71);
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n383), .Q(n15[2]));
    not g155(n78 ,n15[5]);
    nor g156(n559 ,n544 ,n1);
    nor g157(n438 ,n434 ,n436);
    xnor g158(n483 ,n7[0] ,n8[0]);
    nor g159(n181 ,n130 ,n179);
    nor g160(n281 ,n193 ,n195);
    nor g161(n509 ,n168 ,n169);
    nor g162(n399 ,n193 ,n361);
    nor g163(n398 ,n193 ,n353);
    nor g164(n526 ,n118 ,n119);
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n474), .Q(n6[32]));
    nor g166(n113 ,n82 ,n111);
    buf g167(n3[13], n3[15]);
    nor g168(n371 ,n197 ,n279);
    not g169(n75 ,n15[3]);
    not g170(n209 ,n507);
    nor g171(n145 ,n137 ,n142);
    nor g172(n374 ,n232 ,n332);
    not g173(n206 ,n16[47]);
    or g174(n339 ,n299 ,n302);
    nor g175(n415 ,n275 ,n355);
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n553), .Q(n17[4]));
    or g177(n329 ,n249 ,n251);
    not g178(n199 ,n16[63]);
    or g179(n22 ,n15[15] ,n15[14]);
    buf g180(n3[43], n3[47]);
    nor g181(n459 ,n243 ,n455);
    not g182(n219 ,n524);
    nor g183(n21 ,n15[1] ,n15[0]);
    nor g184(n451 ,n406 ,n438);
    not g185(n37 ,n10[9]);
    nor g186(n106 ,n15[7] ,n104);
    or g187(n46 ,n36 ,n35);
    not g188(n303 ,n302);
    nor g189(n278 ,n243 ,n11[1]);
    nor g190(n525 ,n121 ,n122);
    not g191(n230 ,n523);
    not g192(n79 ,n15[8]);
    or g193(n51 ,n37 ,n50);
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n367), .Q(n10[7]));
    not g195(n133 ,n10[2]);
    or g196(n59 ,n15[9] ,n15[8]);
    nor g197(n175 ,n139 ,n173);
    not g198(n131 ,n10[3]);
    not g199(n182 ,n181);
    or g200(n498 ,n479 ,n488);
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n562), .Q(n17[1]));
    not g202(n264 ,n15[4]);
    dff g203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n472), .Q(n6[40]));
    nor g204(n286 ,n226 ,n498);
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n577), .Q(n17[19]));
    nor g206(n563 ,n543 ,n1);
    buf g207(n3[22], n3[23]);
    not g208(n143 ,n10[12]);
    not g209(n82 ,n15[9]);
    not g210(n261 ,n15[6]);
    or g211(n548 ,n17[4] ,n1);
    not g212(n256 ,n15[15]);
    or g213(n42 ,n10[11] ,n10[10]);
    not g214(n208 ,n505);
    not g215(n231 ,n511);
    nor g216(n378 ,n213 ,n332);
    nor g217(n92 ,n77 ,n90);
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n309), .Q(n4[0]));
    or g219(n24 ,n15[9] ,n15[8]);
    buf g220(n3[27], n3[31]);
    xor g221(n358 ,n499 ,n13[0]);
    buf g222(n3[35], n3[39]);
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n308), .Q(n4[1]));
    or g224(n467 ,n459 ,n452);
    nor g225(n364 ,n238 ,n332);
    not g226(n263 ,n15[3]);
    nor g227(n160 ,n129 ,n158);
    not g228(n173 ,n172);
    buf g229(n3[34], n3[39]);
    not g230(n152 ,n151);
    buf g231(n3[3], n3[7]);
    not g232(n265 ,n15[13]);
    nor g233(n379 ,n216 ,n332);
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n468), .Q(n11[1]));
    not g235(n84 ,n15[14]);
    or g236(n475 ,n449 ,n464);
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n282), .Q(n5[7]));
    nor g238(n321 ,n271 ,n194);
    nor g239(n443 ,n16[63] ,n441);
    nor g240(n445 ,n16[47] ,n441);
    or g241(n385 ,n193 ,n362);
    nor g242(n277 ,n245 ,n12[0]);
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n558), .Q(n17[13]));
    buf g244(n3[38], n3[39]);
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n310), .Q(n5[6]));
    not g246(n244 ,n11[1]);
    or g247(n317 ,n247 ,n250);
    nor g248(n118 ,n15[11] ,n116);
    not g249(n546 ,n17[19]);
    not g250(n496 ,n521);
    not g251(n195 ,n16[7]);
    not g252(n216 ,n514);
    or g253(n520 ,n43 ,n54);
    nor g254(n177 ,n10[12] ,n175);
    dff g255(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n473), .Q(n6[0]));
    nor g256(n523 ,n127 ,n128);
    not g257(n234 ,n503);
    not g258(n36 ,n10[8]);
    nor g259(n180 ,n10[13] ,n178);
    nor g260(n183 ,n10[14] ,n181);
    or g261(n69 ,n15[15] ,n67);
    nor g262(n508 ,n165 ,n166);
    or g263(n275 ,n244 ,n11[0]);
    or g264(n31 ,n18 ,n29);
    dff g265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n570), .Q(n16[23]));
    not g266(n232 ,n508);
    nor g267(n432 ,n284 ,n420);
    xor g268(n574 ,n17[5] ,n2[5]);
    nor g269(n533 ,n97 ,n98);
    nor g270(n63 ,n55 ,n58);
    nor g271(n192 ,n187 ,n190);
    buf g272(n3[59], n3[63]);
    nor g273(n504 ,n153 ,n154);
    nor g274(n98 ,n76 ,n96);
    nor g275(n458 ,n244 ,n455);
    not g276(n545 ,n17[18]);
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n551), .Q(n17[11]));
    buf g278(n3[18], n3[23]);
    xnor g279(n566 ,n17[11] ,n17[15]);
    buf g280(n3[42], n3[47]);
    nor g281(n290 ,n214 ,n498);
    nor g282(n125 ,n74 ,n123);
    or g283(n61 ,n15[7] ,n15[6]);
    nor g284(n29 ,n23 ,n28);
    not g285(n210 ,n517);
    buf g286(n3[14], n3[15]);
    dff g287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n571), .Q(n16[15]));
    not g288(n137 ,n10[1]);
    or g289(n577 ,n1 ,n576);
    not g290(n268 ,n5[3]);
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n559), .Q(n17[9]));
    nor g292(n320 ,n270 ,n194);
    buf g293(n3[46], n3[47]);
    buf g294(n3[2], n3[7]);
    nor g295(n529 ,n109 ,n110);
    xnor g296(n423 ,n362 ,n12[0]);
    buf g297(n3[16], n3[23]);
    not g298(n93 ,n92);
    nor g299(n151 ,n131 ,n149);
    nor g300(n313 ,n259 ,n194);
    nor g301(n295 ,n230 ,n498);
    nor g302(n391 ,n242 ,n356);
    nor g303(n524 ,n124 ,n125);
    nor g304(n530 ,n106 ,n107);
    not g305(n213 ,n513);
    not g306(n253 ,n5[4]);
    nor g307(n124 ,n15[13] ,n122);
    or g308(n516 ,n69 ,n72);
    nor g309(n561 ,n542 ,n1);
    nor g310(n389 ,n193 ,n343);
    not g311(n130 ,n10[13]);
    not g312(n141 ,n10[10]);
    nor g313(n283 ,n235 ,n498);
    nor g314(n308 ,n247 ,n193);
    nor g315(n400 ,n277 ,n359);
    nor g316(n412 ,n210 ,n361);
    nor g317(n454 ,n193 ,n439);
    nor g318(n463 ,n200 ,n453);
    nor g319(n305 ,n268 ,n193);
    not g320(n224 ,n512);
    dff g321(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n548), .Q(n17[3]));
    nor g322(n421 ,n410 ,n412);
    nor g323(n171 ,n10[10] ,n169);
    buf g324(n3[10], n3[15]);
    not g325(n140 ,n10[14]);
    xor g326(n491 ,n489 ,n490);
    not g327(n18 ,n15[6]);
    nor g328(n348 ,n322 ,n286);
    nor g329(n535 ,n91 ,n92);
    not g330(n406 ,n405);
    not g331(n197 ,n2[0]);
    nor g332(n457 ,n195 ,n453);
    not g333(n240 ,n518);
    nor g334(n469 ,n450 ,n456);
    or g335(n547 ,n17[13] ,n1);
    or g336(n27 ,n22 ,n26);
    nor g337(n95 ,n75 ,n93);
    nor g338(n352 ,n324 ,n290);
    not g339(n271 ,n15[10]);
    nor g340(n449 ,n16[15] ,n441);
    not g341(n80 ,n15[7]);
    nor g342(n456 ,n301 ,n454);
    not g343(n164 ,n163);
    nor g344(n511 ,n174 ,n175);
    dff g345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n392), .Q(n15[10]));
    nor g346(n331 ,n265 ,n194);
    nor g347(n354 ,n10[0] ,n332);
    or g348(n340 ,n274 ,n276);
    nor g349(n433 ,n193 ,n423);
    xnor g350(n3[39] ,n491 ,n6[32]);
    not g351(n76 ,n15[4]);
    not g352(n227 ,n509);
    or g353(n500 ,n495 ,n492);
    xor g354(n334 ,n498 ,n15[0]);
    nor g355(n404 ,n193 ,n345);
    dff g356(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n433), .Q(n12[0]));
    not g357(n222 ,n506);
    xnor g358(n486 ,n481 ,n480);
    nor g359(n347 ,n313 ,n294);
    not g360(n81 ,n15[1]);
    nor g361(n392 ,n193 ,n360);
    dff g362(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n549), .Q(n17[8]));
    not g363(n250 ,n4[2]);
    buf g364(n3[28], n3[31]);
    dff g365(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n547), .Q(n17[12]));
    dff g366(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n568), .Q(n16[39]));
    nor g367(n373 ,n234 ,n332);
    nor g368(n396 ,n193 ,n351);
    nor g369(n556 ,n537 ,n1);
    nor g370(n47 ,n10[1] ,n44);
    nor g371(n409 ,n249 ,n362);
    nor g372(n519 ,n189 ,n188);
    nor g373(n68 ,n15[2] ,n65);
    nor g374(n103 ,n15[6] ,n101);
    dff g375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n304), .Q(n5[5]));
    not g376(n242 ,n11[0]);
    nor g377(n319 ,n263 ,n194);
    not g378(n241 ,n533);
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n372), .Q(n10[4]));
    nor g380(n417 ,n415 ,n402);
    nor g381(n401 ,n193 ,n334);
    nor g382(n338 ,n11[2] ,n299);
    nor g383(n318 ,n254 ,n194);
    buf g384(n3[12], n3[15]);
    nor g385(n447 ,n16[31] ,n441);
    or g386(n474 ,n446 ,n463);
    nor g387(n153 ,n10[4] ,n151);
    not g388(n56 ,n15[4]);
    buf g389(n3[29], n3[31]);
    not g390(n196 ,n8[1]);
    nor g391(n503 ,n150 ,n151);
    buf g392(n3[19], n3[23]);
    not g393(n73 ,n15[6]);
    nor g394(n280 ,n245 ,n193);
    dff g395(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n280), .Q(n7[0]));
    xor g396(n576 ,n566 ,n567);
    nor g397(n276 ,n244 ,n516);
    nor g398(n534 ,n94 ,n95);
    xor g399(n569 ,n17[3] ,n2[3]);
    xnor g400(n3[31] ,n491 ,n6[24]);
    not g401(n58 ,n15[0]);
    not g402(n269 ,n15[14]);
    xor g403(n570 ,n17[2] ,n2[2]);
    not g404(n361 ,n362);
    buf g405(n3[58], n3[63]);
    not g406(n494 ,n5[5]);
    nor g407(n316 ,n269 ,n194);
    nor g408(n166 ,n135 ,n164);
    nor g409(n273 ,n8[0] ,n11[0]);
    dff g410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n388), .Q(n15[14]));
    nor g411(n147 ,n10[2] ,n145);
    nor g412(n431 ,n193 ,n421);
    buf g413(n3[25], n3[31]);
    xor g414(n568 ,n17[4] ,n2[4]);
    nor g415(n558 ,n540 ,n1);
    dff g416(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n364), .Q(n10[1]));
    or g417(n473 ,n448 ,n457);
    nor g418(n312 ,n198 ,n194);
    xor g419(n515 ,n10[15] ,n184);
    dff g420(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n384), .Q(n15[1]));
    not g421(n212 ,n515);
    or g422(n422 ,n299 ,n391);
    not g423(n540 ,n17[14]);
    nor g424(n91 ,n15[2] ,n89);
    nor g425(n464 ,n202 ,n453);
    nor g426(n88 ,n15[1] ,n15[0]);
    not g427(n99 ,n98);
    not g428(n167 ,n166);
    nor g429(n390 ,n193 ,n344);
    nor g430(n403 ,n193 ,n358);
    not g431(n238 ,n501);
    or g432(n30 ,n25 ,n27);
    not g433(n74 ,n15[13]);
    not g434(n142 ,n10[0]);
    nor g435(n383 ,n193 ,n336);
    not g436(n228 ,n531);
    not g437(n226 ,n529);
    nor g438(n387 ,n193 ,n341);
    nor g439(n297 ,n221 ,n498);
    not g440(n258 ,n15[5]);
    nor g441(n536 ,n89 ,n88);
    not g442(n205 ,n15[2]);
    not g443(n132 ,n10[4]);
    dff g444(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n574), .Q(n16[47]));
    dff g445(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n396), .Q(n15[6]));
    nor g446(n122 ,n87 ,n120);
    nor g447(n307 ,n266 ,n193);
    dff g448(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n550), .Q(n17[7]));
    nor g449(n375 ,n231 ,n332);
    dff g450(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n563), .Q(n17[5]));
    nor g451(n342 ,n316 ,n295);
    not g452(n139 ,n10[11]);
    or g453(n471 ,n444 ,n461);
    not g454(n266 ,n4[1]);
    nor g455(n288 ,n211 ,n498);
    nor g456(n121 ,n15[12] ,n119);
    xor g457(n575 ,n17[6] ,n2[6]);
    nor g458(n397 ,n193 ,n352);
    xor g459(n573 ,n17[7] ,n2[7]);
    nor g460(n450 ,n11[0] ,n439);
    dff g461(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n306), .Q(n5[3]));
    not g462(n176 ,n175);
    not g463(n102 ,n101);
    nor g464(n376 ,n224 ,n332);
    not g465(n96 ,n95);
    nor g466(n346 ,n212 ,n332);
    nor g467(n461 ,n204 ,n453);
    not g468(n155 ,n154);
    buf g469(n3[4], n3[7]);
    dff g470(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n569), .Q(n16[31]));
    or g471(n279 ,n245 ,n8[1]);
    nor g472(n408 ,n252 ,n362);
    nor g473(n326 ,n243 ,n197);
    buf g474(n3[11], n3[15]);
    or g475(n43 ,n10[15] ,n10[14]);
    not g476(n77 ,n15[2]);
    not g477(n19 ,n15[2]);
    nor g478(n94 ,n15[3] ,n92);
    not g479(n38 ,n10[3]);
    nor g480(n337 ,n312 ,n283);
    nor g481(n363 ,n223 ,n332);
    buf g482(n3[48], n3[55]);
    nor g483(n394 ,n193 ,n348);
    nor g484(n178 ,n143 ,n176);
    nor g485(n414 ,n239 ,n361);
    nor g486(n345 ,n320 ,n288);
    not g487(n233 ,n510);
    not g488(n542 ,n17[11]);
    or g489(n355 ,n500 ,n317);
    not g490(n179 ,n178);
    buf g491(n3[1], n3[7]);
    nor g492(n154 ,n132 ,n152);
    nor g493(n446 ,n16[39] ,n441);
    nor g494(n299 ,n242 ,n244);
    nor g495(n272 ,n8[0] ,n499);
    nor g496(n188 ,n12[1] ,n12[0]);
    or g497(n499 ,n478 ,n498);
    dff g498(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n404), .Q(n15[11]));
    or g499(n551 ,n17[12] ,n1);
    nor g500(n49 ,n38 ,n47);
    not g501(n136 ,n10[7]);
    dff g502(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n397), .Q(n15[5]));
    xor g503(n490 ,n499 ,n483);
    or g504(n420 ,n260 ,n400);
    buf g505(n3[9], n3[15]);
    not g506(n85 ,n15[10]);
    dff g507(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n430), .Q(n12[2]));
    nor g508(n460 ,n199 ,n453);
    nor g509(n311 ,n205 ,n194);
    nor g510(n349 ,n314 ,n285);
    xnor g511(n3[47] ,n491 ,n6[40]);
    or g512(n437 ,n193 ,n432);
    nor g513(n322 ,n262 ,n194);
    nor g514(n293 ,n225 ,n498);
    not g515(n138 ,n10[9]);
    buf g516(n3[54], n3[55]);
    dff g517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n301), .Q(n8[0]));
    buf g518(n3[36], n3[39]);
    or g519(n34 ,n15[7] ,n33);
    nor g520(n505 ,n156 ,n157);
    dff g521(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n564), .Q(n17[18]));
    xnor g522(n3[63] ,n491 ,n6[56]);
    or g523(n25 ,n15[13] ,n15[12]);
    or g524(n468 ,n458 ,n451);
    xnor g525(n480 ,n13[0] ,n14[0]);
    or g526(n52 ,n46 ,n51);
    nor g527(n425 ,n338 ,n385);
    buf g528(n3[37], n3[39]);
    dff g529(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n377), .Q(n10[10]));
    not g530(n187 ,n12[2]);
    dff g531(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n399), .Q(n8[3]));
    dff g532(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n565), .Q(n17[14]));
    not g533(n185 ,n12[1]);
    or g534(n436 ,n435 ,n427);
    not g535(n170 ,n169);
    not g536(n539 ,n17[2]);
    nor g537(n335 ,n319 ,n297);
    dff g538(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n469), .Q(n11[0]));
    or g539(n488 ,n5[6] ,n487);
    dff g540(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n398), .Q(n15[4]));
    dff g541(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n573), .Q(n16[63]));
    dff g542(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n557), .Q(n17[17]));
    nor g543(n189 ,n185 ,n186);
    dff g544(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n555), .Q(n17[0]));
    nor g545(n298 ,n217 ,n498);
    not g546(n229 ,n2[1]);
    not g547(n235 ,n536);
    not g548(n217 ,n525);
    not g549(n300 ,n299);
    buf g550(n3[33], n3[39]);
    nor g551(n172 ,n141 ,n170);
    buf g552(n3[51], n3[55]);
    not g553(n441 ,n440);
    or g554(n66 ,n59 ,n61);
    not g555(n149 ,n148);
    dff g556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n470), .Q(n6[56]));
    nor g557(n434 ,n407 ,n422);
    nor g558(n148 ,n133 ,n146);
    not g559(n202 ,n16[15]);
    not g560(n245 ,n8[0]);
    not g561(n198 ,n15[1]);
    nor g562(n116 ,n85 ,n114);
    or g563(n33 ,n30 ,n32);
    nor g564(n512 ,n177 ,n178);
    dff g565(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n393), .Q(n15[9]));
    not g566(n493 ,n5[7]);
    nor g567(n440 ,n437 ,n428);
    nor g568(n393 ,n193 ,n347);
    nor g569(n325 ,n264 ,n194);
    nor g570(n502 ,n147 ,n148);
    nor g571(n386 ,n193 ,n333);
    or g572(n428 ,n8[3] ,n424);
    nor g573(n165 ,n10[8] ,n163);
    dff g574(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n556), .Q(n17[6]));
    not g575(n247 ,n4[0]);
    nor g576(n327 ,n248 ,n245);
    not g577(n220 ,n527);
    buf g578(n3[40], n3[47]);
    not g579(n55 ,n15[1]);
    nor g580(n284 ,n247 ,n8[1]);
    buf g581(n3[56], n3[63]);
    dff g582(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n354), .Q(n10[0]));
    buf g583(n3[24], n3[31]);
    dff g584(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n382), .Q(n15[3]));
    nor g585(n444 ,n16[55] ,n441);
    nor g586(n287 ,n220 ,n498);
    or g587(n67 ,n60 ,n62);
    nor g588(n452 ,n426 ,n438);
    nor g589(n89 ,n81 ,n86);
    not g590(n207 ,n530);
    or g591(n54 ,n48 ,n53);
    xnor g592(n489 ,n486 ,n482);
    nor g593(n128 ,n84 ,n126);
    buf g594(n3[45], n3[47]);
    or g595(n45 ,n39 ,n40);
    not g596(n129 ,n10[6]);
    not g597(n478 ,n516);
    nor g598(n429 ,n193 ,n416);
    buf g599(n3[57], n3[63]);
    nor g600(n159 ,n10[6] ,n157);
    buf g601(n3[52], n3[55]);
    nor g602(n169 ,n138 ,n167);
    or g603(n44 ,n10[2] ,n10[0]);
    not g604(n126 ,n125);
    nor g605(n285 ,n207 ,n498);
    nor g606(n163 ,n136 ,n161);
    nor g607(n507 ,n162 ,n163);
    not g608(n215 ,n504);
    buf g609(n3[44], n3[47]);
    not g610(n495 ,n4[1]);
    or g611(n485 ,n493 ,n484);
    not g612(n439 ,n438);
    xor g613(n571 ,n17[1] ,n2[1]);
    dff g614(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n575), .Q(n16[55]));
    xor g615(n522 ,n15[15] ,n128);
    nor g616(n427 ,n11[2] ,n417);
    or g617(n330 ,n236 ,n229);
    not g618(n270 ,n15[11]);
    or g619(n550 ,n17[8] ,n1);
    nor g620(n353 ,n325 ,n296);
    nor g621(n150 ,n10[3] ,n148);
    nor g622(n532 ,n100 ,n101);
    or g623(n407 ,n243 ,n340);
    nor g624(n343 ,n331 ,n292);
    not g625(n543 ,n17[6]);
    nor g626(n168 ,n10[9] ,n166);
    not g627(n111 ,n110);
    dff g628(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n374), .Q(n10[8]));
    nor g629(n50 ,n10[4] ,n49);
    or g630(n521 ,n24 ,n34);
    nor g631(n310 ,n267 ,n193);
    nor g632(n430 ,n193 ,n418);
    or g633(n555 ,n17[1] ,n1);
    nor g634(n53 ,n45 ,n52);
    dff g635(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n376), .Q(n10[12]));
    buf g636(n3[32], n3[39]);
    nor g637(n410 ,n251 ,n362);
    nor g638(n557 ,n545 ,n1);
    dff g639(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n395), .Q(n15[7]));
    nor g640(n506 ,n159 ,n160);
    dff g641(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n560), .Q(n17[2]));
    nor g642(n367 ,n209 ,n332);
    buf g643(n3[26], n3[31]);
    or g644(n64 ,n57 ,n56);
    or g645(n71 ,n66 ,n70);
    nor g646(n289 ,n228 ,n498);
    not g647(n105 ,n104);
    not g648(n194 ,n498);
    dff g649(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n373), .Q(n10[3]));
    or g650(n381 ,n8[2] ,n371);
    dff g651(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n475), .Q(n6[8]));
    nor g652(n274 ,n194 ,n11[0]);
    nor g653(n109 ,n15[8] ,n107);
    nor g654(n513 ,n180 ,n181);
    nor g655(n368 ,n222 ,n332);
    not g656(n260 ,n8[2]);
    nor g657(n304 ,n253 ,n193);
    not g658(n214 ,n532);
    dff g659(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n375), .Q(n10[11]));
    nor g660(n315 ,n256 ,n194);
    xnor g661(n482 ,n9[0] ,n10[0]);
    not g662(n254 ,n15[12]);
    dff g663(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n378), .Q(n10[13]));
    not g664(n537 ,n17[7]);
    buf g665(n3[60], n3[63]);
    or g666(n549 ,n17[9] ,n1);
    or g667(n476 ,n442 ,n465);
    buf g668(n3[6], n3[7]);
    nor g669(n411 ,n196 ,n350);
    buf g670(n3[50], n3[55]);
    or g671(n62 ,n15[11] ,n15[10]);
    nor g672(n395 ,n193 ,n349);
    dff g673(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n368), .Q(n10[6]));
    or g674(n402 ,n369 ,n370);
    not g675(n211 ,n526);
    nor g676(n104 ,n73 ,n102);
    not g677(n426 ,n425);
    not g678(n193 ,n1);
    or g679(n552 ,n17[17] ,n1);
    or g680(n487 ,n4[2] ,n485);
    nor g681(n292 ,n219 ,n498);
    not g682(n20 ,n15[5]);
    nor g683(n442 ,n16[23] ,n441);
    nor g684(n514 ,n183 ,n184);
    nor g685(n97 ,n15[4] ,n95);
    dff g686(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n429), .Q(n12[1]));
    nor g687(n100 ,n15[5] ,n98);
    not g688(n541 ,n17[3]);
    not g689(n249 ,n12[2]);
    buf g690(n3[17], n3[23]);
    not g691(n123 ,n122);
    nor g692(n282 ,n257 ,n193);
    nor g693(n527 ,n115 ,n116);
    nor g694(n362 ,n243 ,n300);
    dff g695(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n390), .Q(n15[12]));
    not g696(n225 ,n522);
    dff g697(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n403), .Q(n13[0]));
    not g698(n190 ,n189);
    nor g699(n560 ,n541 ,n1);
    nor g700(n418 ,n409 ,n413);
    nor g701(n382 ,n193 ,n335);
    nor g702(n291 ,n237 ,n498);
    or g703(n479 ,n494 ,n5[4]);
    not g704(n83 ,n15[11]);
    not g705(n223 ,n502);
    nor g706(n341 ,n315 ,n293);
    nor g707(n127 ,n15[14] ,n125);
    not g708(n455 ,n454);
    not g709(n221 ,n534);
    nor g710(n531 ,n103 ,n104);
    xnor g711(n3[23] ,n491 ,n6[16]);
    xnor g712(n3[55] ,n491 ,n6[48]);
    nor g713(n356 ,n328 ,n329);
    nor g714(n370 ,n496 ,n303);
endmodule
