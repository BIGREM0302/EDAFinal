module top(n0, n1, n2, n3, n5, n8, n6, n9, n4, n7, n10, n11, n12, n13);
    input n0, n1;
    input [15:0] n2;
    input [7:0] n3, n4;
    input [3:0] n5, n6, n7;
    input [5:0] n8;
    input [1:0] n9;
    output [7:0] n10;
    output [3:0] n11;
    output [1:0] n12;
    output n13;
    wire n0, n1;
    wire [15:0] n2;
    wire [7:0] n3, n4;
    wire [3:0] n5, n6, n7;
    wire [5:0] n8;
    wire [1:0] n9;
    wire [7:0] n10;
    wire [3:0] n11;
    wire [1:0] n12;
    wire n13;
    wire [15:0] n14;
    wire [7:0] n15;
    wire [7:0] n16;
    wire [7:0] n17;
    wire [7:0] n18;
    wire [15:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [7:0] n22;
    wire [15:0] n23;
    wire [7:0] n24;
    wire [15:0] n25;
    wire [15:0] n26;
    wire [15:0] n27;
    wire [15:0] n28;
    wire [15:0] n29;
    wire [15:0] n30;
    wire [7:0] n31;
    wire [7:0] n32;
    wire [7:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [7:0] n36;
    wire [2:0] n37;
    wire [2:0] n38;
    wire [7:0] n39;
    wire [7:0] n40;
    wire [7:0] n41;
    wire [7:0] n42;
    wire [7:0] n43;
    wire [7:0] n44;
    wire [7:0] n45;
    wire [7:0] n46;
    wire [7:0] n47;
    wire n48, n49, n50, n51, n52, n53, n54, n55;
    wire n56, n57, n58, n59, n60, n61, n62, n63;
    wire n64, n65, n66, n67, n68, n69, n70, n71;
    wire n72, n73, n74, n75, n76, n77, n78, n79;
    wire n80, n81, n82, n83, n84, n85, n86, n87;
    wire n88, n89, n90, n91, n92, n93, n94, n95;
    wire n96, n97, n98, n99, n100, n101, n102, n103;
    wire n104, n105, n106, n107, n108, n109, n110, n111;
    wire n112, n113, n114, n115, n116, n117, n118, n119;
    wire n120, n121, n122, n123, n124, n125, n126, n127;
    wire n128, n129, n130, n131, n132, n133, n134, n135;
    wire n136, n137, n138, n139, n140, n141, n142, n143;
    wire n144, n145, n146, n147, n148, n149, n150, n151;
    wire n152, n153, n154, n155, n156, n157, n158, n159;
    wire n160, n161, n162, n163, n164, n165, n166, n167;
    wire n168, n169, n170, n171, n172, n173, n174, n175;
    wire n176, n177, n178, n179, n180, n181, n182, n183;
    wire n184, n185, n186, n187, n188, n189, n190, n191;
    wire n192, n193, n194, n195, n196, n197, n198, n199;
    wire n200, n201, n202, n203, n204, n205, n206, n207;
    wire n208, n209, n210, n211, n212, n213, n214, n215;
    wire n216, n217, n218, n219, n220, n221, n222, n223;
    wire n224, n225, n226, n227, n228, n229, n230, n231;
    wire n232, n233, n234, n235, n236, n237, n238, n239;
    wire n240, n241, n242, n243, n244, n245, n246, n247;
    wire n248, n249, n250, n251, n252, n253, n254, n255;
    wire n256, n257, n258, n259, n260, n261, n262, n263;
    wire n264, n265, n266, n267, n268, n269, n270, n271;
    wire n272, n273, n274, n275, n276, n277, n278, n279;
    wire n280, n281, n282, n283, n284, n285, n286, n287;
    wire n288, n289, n290, n291, n292, n293, n294, n295;
    wire n296, n297, n298, n299, n300, n301, n302, n303;
    wire n304, n305, n306, n307, n308, n309, n310, n311;
    wire n312, n313, n314, n315, n316, n317, n318, n319;
    wire n320, n321, n322, n323, n324, n325, n326, n327;
    wire n328, n329, n330, n331, n332, n333, n334, n335;
    wire n336, n337, n338, n339, n340, n341, n342, n343;
    wire n344, n345, n346, n347, n348, n349, n350, n351;
    wire n352, n353, n354, n355, n356, n357, n358, n359;
    wire n360, n361, n362, n363, n364, n365, n366, n367;
    wire n368, n369, n370, n371, n372, n373, n374, n375;
    wire n376, n377, n378, n379, n380, n381, n382, n383;
    wire n384, n385, n386, n387, n388, n389, n390, n391;
    wire n392, n393, n394, n395, n396, n397, n398, n399;
    wire n400, n401, n402, n403, n404, n405, n406, n407;
    wire n408, n409, n410, n411, n412, n413, n414, n415;
    wire n416, n417, n418, n419, n420, n421, n422, n423;
    wire n424, n425, n426, n427, n428, n429, n430, n431;
    wire n432, n433, n434, n435, n436, n437, n438, n439;
    wire n440, n441, n442, n443, n444, n445, n446, n447;
    wire n448, n449, n450, n451, n452, n453, n454, n455;
    wire n456, n457, n458, n459, n460, n461, n462, n463;
    wire n464, n465, n466, n467, n468, n469, n470, n471;
    wire n472, n473, n474, n475, n476, n477, n478, n479;
    wire n480, n481, n482, n483, n484, n485, n486, n487;
    wire n488, n489, n490, n491, n492, n493, n494, n495;
    wire n496, n497, n498, n499, n500, n501, n502, n503;
    wire n504, n505, n506, n507, n508, n509, n510, n511;
    wire n512, n513, n514, n515, n516, n517, n518, n519;
    wire n520, n521, n522, n523, n524, n525, n526, n527;
    wire n528, n529, n530, n531, n532, n533, n534, n535;
    xor g0(n147 ,n40[3] ,n6[1]);
    xor g1(n133 ,n2[4] ,n3[4]);
    not g2(n451 ,n17[7]);
    nor g3(n290 ,n195 ,n210);
    nor g4(n274 ,n453 ,n215);
    dff g5(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[7]), .Q(n24[7]));
    not g6(n52 ,n30[5]);
    or g7(n346 ,n323 ,n319);
    nor g8(n350 ,n338 ,n336);
    nor g9(n240 ,n462 ,n212);
    not g10(n495 ,n350);
    xor g11(n148 ,n27[3] ,n42[3]);
    xnor g12(n160 ,n5[0] ,n111);
    or g13(n303 ,n293 ,n273);
    xor g14(n95 ,n39[3] ,n6[0]);
    xnor g15(n391 ,n30[0] ,n380);
    not g16(n491 ,n15[2]);
    xor g17(n94 ,n34[4] ,n8[4]);
    or g18(n421 ,n213 ,n417);
    nor g19(n262 ,n454 ,n209);
    xnor g20(n159 ,n9[0] ,n71);
    not g21(n193 ,n36[1]);
    nor g22(n272 ,n451 ,n210);
    or g23(n529 ,n525 ,n524);
    not g24(n462 ,n23[2]);
    nor g25(n286 ,n450 ,n209);
    or g26(n341 ,n329 ,n315);
    dff g27(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[1]), .Q(n19[1]));
    not g28(n58 ,n30[7]);
    xnor g29(n379 ,n375 ,n33[2]);
    not g30(n457 ,n24[3]);
    xor g31(n83 ,n43[2] ,n7[0]);
    dff g32(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[5]), .Q(n23[7]));
    dff g33(.RN(n1), .SN(1'b1), .CK(n0), .D(n169), .Q(n34[3]));
    or g34(n66 ,n58 ,n30[6]);
    dff g35(.RN(n1), .SN(1'b1), .CK(n0), .D(n130), .Q(n20[2]));
    dff g36(.RN(n1), .SN(1'b1), .CK(n0), .D(n136), .Q(n36[0]));
    not g37(n56 ,n30[3]);
    dff g38(.RN(n1), .SN(1'b1), .CK(n0), .D(n126), .Q(n18[1]));
    not g39(n471 ,n14[3]);
    xnor g40(n387 ,n32[2] ,n379);
    or g41(n299 ,n228 ,n262);
    nor g42(n247 ,n471 ,n214);
    or g43(n505 ,n340 ,n428);
    dff g44(.RN(n1), .SN(1'b1), .CK(n0), .D(n157), .Q(n26[0]));
    dff g45(.RN(n1), .SN(1'b1), .CK(n0), .D(n493), .Q(n10[4]));
    xnor g46(n175 ,n120 ,n32[2]);
    or g47(n318 ,n284 ,n283);
    dff g48(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[4]), .Q(n29[6]));
    xnor g49(n157 ,n8[4] ,n73);
    xor g50(n139 ,n29[1] ,n41[1]);
    or g51(n330 ,n285 ,n281);
    dff g52(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[2]), .Q(n29[4]));
    or g53(n308 ,n234 ,n233);
    not g54(n184 ,n36[0]);
    dff g55(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[11]), .Q(n25[1]));
    or g56(n149 ,n65 ,n61);
    xor g57(n127 ,n46[3] ,n4[7]);
    nor g58(n219 ,n429 ,n208);
    xor g59(n98 ,n39[1] ,n4[0]);
    or g60(n295 ,n243 ,n238);
    xnor g61(n73 ,n2[8] ,n3[4]);
    dff g62(.RN(n1), .SN(1'b1), .CK(n0), .D(n140), .Q(n30[6]));
    dff g63(.RN(n1), .SN(1'b1), .CK(n0), .D(n164), .Q(n36[3]));
    nor g64(n254 ,n475 ,n212);
    dff g65(.RN(n1), .SN(1'b1), .CK(n0), .D(n174), .Q(n28[0]));
    or g66(n422 ,n213 ,n419);
    dff g67(.RN(n1), .SN(1'b1), .CK(n0), .D(n176), .Q(n32[3]));
    not g68(n453 ,n25[2]);
    nor g69(n217 ,n487 ,n208);
    nor g70(n233 ,n465 ,n212);
    dff g71(.RN(n1), .SN(1'b1), .CK(n0), .D(n129), .Q(n20[3]));
    dff g72(.RN(n1), .SN(1'b1), .CK(n0), .D(n499), .Q(n10[2]));
    or g73(n339 ,n300 ,n298);
    nor g74(n242 ,n445 ,n213);
    nor g75(n230 ,n490 ,n212);
    nor g76(n279 ,n437 ,n216);
    not g77(n436 ,n29[7]);
    not g78(n180 ,n37[1]);
    not g79(n480 ,n20[2]);
    or g80(n154 ,n67 ,n152);
    xor g81(n362 ,n498 ,n36[1]);
    nor g82(n418 ,n293 ,n413);
    dff g83(.RN(n1), .SN(1'b1), .CK(n0), .D(n153), .Q(n17[2]));
    nor g84(n293 ,n440 ,n213);
    nor g85(n280 ,n457 ,n209);
    dff g86(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[3]), .Q(n28[5]));
    nor g87(n253 ,n192 ,n214);
    not g88(n60 ,n30[14]);
    xor g89(n110 ,n41[1] ,n7[2]);
    xnor g90(n367 ,n359 ,n35[2]);
    not g91(n55 ,n30[1]);
    dff g92(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[3]), .Q(n28[1]));
    or g93(n326 ,n291 ,n224);
    or g94(n68 ,n55 ,n30[0]);
    nor g95(n224 ,n486 ,n208);
    dff g96(.RN(n1), .SN(1'b1), .CK(n0), .D(n143), .Q(n35[1]));
    nor g97(n419 ,n294 ,n414);
    dff g98(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[6]), .Q(n22[6]));
    not g99(n192 ,n35[3]);
    dff g100(.RN(n1), .SN(1'b1), .CK(n0), .D(n148), .Q(n21[3]));
    nor g101(n277 ,n438 ,n216);
    or g102(n322 ,n288 ,n287);
    nor g103(n535 ,n534 ,n533);
    dff g104(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[6]), .Q(n17[6]));
    not g105(n472 ,n14[6]);
    xnor g106(n118 ,n5[2] ,n8[2]);
    or g107(n405 ,n213 ,n397);
    xnor g108(n124 ,n5[2] ,n36[2]);
    xnor g109(n404 ,n388 ,n31[3]);
    xor g110(n78 ,n46[2] ,n7[3]);
    xnor g111(n113 ,n2[2] ,n3[2]);
    dff g112(.RN(n1), .SN(1'b1), .CK(n0), .D(n134), .Q(n18[2]));
    dff g113(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[4]), .Q(n27[6]));
    not g114(n446 ,n26[2]);
    or g115(n399 ,n241 ,n396);
    dff g116(.RN(n1), .SN(1'b1), .CK(n0), .D(n168), .Q(n34[2]));
    nor g117(n275 ,n431 ,n216);
    nor g118(n51 ,n49 ,n48);
    or g119(n524 ,n519 ,n518);
    dff g120(.RN(n512), .SN(1'b1), .CK(n0), .D(n505), .Q(n47[3]));
    xnor g121(n74 ,n8[2] ,n34[2]);
    not g122(n432 ,n18[2]);
    not g123(n182 ,n32[2]);
    xnor g124(n161 ,n5[3] ,n114);
    dff g125(.RN(n1), .SN(1'b1), .CK(n0), .D(n171), .Q(n19[0]));
    dff g126(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[13]), .Q(n23[1]));
    nor g127(n410 ,n402 ,n406);
    dff g128(.RN(n1), .SN(1'b1), .CK(n0), .D(n14[3]), .Q(n14[5]));
    not g129(n460 ,n18[6]);
    dff g130(.RN(n512), .SN(1'b1), .CK(n0), .D(n508), .Q(n47[0]));
    not g131(n434 ,n29[6]);
    xnor g132(n403 ,n387 ,n31[2]);
    not g133(n414 ,n413);
    xor g134(n126 ,n28[1] ,n40[1]);
    nor g135(n383 ,n216 ,n379);
    not g136(n438 ,n28[7]);
    nor g137(n288 ,n455 ,n215);
    nor g138(n270 ,n186 ,n215);
    not g139(n447 ,n18[7]);
    xor g140(n145 ,n27[1] ,n42[1]);
    xor g141(n136 ,n36[0] ,n5[0]);
    nor g142(n401 ,n189 ,n392);
    xnor g143(n380 ,n378 ,n33[0]);
    dff g144(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[5]), .Q(n29[7]));
    nor g145(n234 ,n472 ,n214);
    or g146(n201 ,n179 ,n37[1]);
    not g147(n448 ,n26[3]);
    nor g148(n223 ,n479 ,n208);
    or g149(n506 ,n335 ,n427);
    nor g150(n398 ,n27[1] ,n389);
    xor g151(n140 ,n2[6] ,n3[6]);
    not g152(n440 ,n27[2]);
    nor g153(n397 ,n27[0] ,n391);
    xor g154(n77 ,n33[2] ,n6[2]);
    dff g155(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[2]), .Q(n30[10]));
    dff g156(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[0]), .Q(n23[2]));
    not g157(n474 ,n22[6]);
    nor g158(n408 ,n209 ,n404);
    xnor g159(n368 ,n360 ,n35[0]);
    dff g160(.RN(n1), .SN(1'b1), .CK(n0), .D(n172), .Q(n27[0]));
    or g161(n333 ,n312 ,n301);
    dff g162(.RN(n512), .SN(1'b1), .CK(n0), .D(n506), .Q(n47[2]));
    not g163(n179 ,n37[2]);
    xnor g164(n375 ,n34[2] ,n367);
    dff g165(.RN(n1), .SN(1'b1), .CK(n0), .D(n81), .Q(n44[3]));
    dff g166(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[7]), .Q(n18[7]));
    xor g167(n359 ,n499 ,n36[2]);
    dff g168(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[5]), .Q(n30[13]));
    not g169(n450 ,n24[1]);
    dff g170(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[6]), .Q(n18[6]));
    or g171(n325 ,n292 ,n290);
    or g172(n215 ,n178 ,n201);
    nor g173(n353 ,n208 ,n351);
    not g174(n486 ,n20[7]);
    dff g175(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[7]), .Q(n22[7]));
    not g176(n459 ,n16[6]);
    dff g177(.RN(n1), .SN(1'b1), .CK(n0), .D(n82), .Q(n44[2]));
    dff g178(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[2]), .Q(n19[4]));
    or g179(n340 ,n328 ,n325);
    xor g180(n89 ,n26[3] ,n43[3]);
    or g181(n310 ,n271 ,n268);
    or g182(n306 ,n226 ,n254);
    or g183(n508 ,n399 ,n415);
    not g184(n454 ,n24[2]);
    nor g185(n199 ,n37[2] ,n37[1]);
    xor g186(n176 ,n32[3] ,n166);
    dff g187(.RN(n1), .SN(1'b1), .CK(n0), .D(n500), .Q(n10[3]));
    nor g188(n50 ,n38[1] ,n38[0]);
    xor g189(n137 ,n28[3] ,n40[3]);
    dff g190(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[6]), .Q(n30[14]));
    or g191(n528 ,n503 ,n505);
    dff g192(.RN(n1), .SN(1'b1), .CK(n0), .D(n87), .Q(n41[3]));
    dff g193(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[2]), .Q(n28[4]));
    or g194(n214 ,n180 ,n203);
    or g195(n334 ,n308 ,n305);
    dff g196(.RN(n1), .SN(1'b1), .CK(n0), .D(n107), .Q(n34[0]));
    dff g197(.RN(n1), .SN(1'b1), .CK(n0), .D(n38[1]), .Q(n37[1]));
    dff g198(.RN(n512), .SN(1'b1), .CK(n0), .D(n501), .Q(n47[7]));
    nor g199(n260 ,n463 ,n209);
    nor g200(n510 ,n51 ,n50);
    or g201(n348 ,n327 ,n322);
    or g202(n393 ,n371 ,n383);
    dff g203(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[5]), .Q(n29[1]));
    dff g204(.RN(n1), .SN(1'b1), .CK(n0), .D(n142), .Q(n30[7]));
    dff g205(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[2]), .Q(n23[4]));
    dff g206(.RN(n1), .SN(1'b1), .CK(n0), .D(n38[2]), .Q(n37[2]));
    nor g207(n372 ,n208 ,n368);
    buf g208(n12[1], 1'b0);
    or g209(n314 ,n279 ,n218);
    dff g210(.RN(n1), .SN(1'b1), .CK(n0), .D(n127), .Q(n46[3]));
    dff g211(.RN(n1), .SN(1'b1), .CK(n0), .D(n109), .Q(n22[2]));
    xor g212(n174 ,n116 ,n117);
    not g213(n518 ,n47[7]);
    xor g214(n360 ,n497 ,n36[0]);
    or g215(n363 ,n211 ,n355);
    or g216(n212 ,n180 ,n202);
    not g217(n469 ,n14[2]);
    dff g218(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[6]), .Q(n20[6]));
    xnor g219(n115 ,n5[0] ,n8[0]);
    xnor g220(n72 ,n2[10] ,n3[5]);
    xor g221(n82 ,n44[2] ,n7[1]);
    dff g222(.RN(n1), .SN(1'b1), .CK(n0), .D(n163), .Q(n30[1]));
    xnor g223(n122 ,n5[3] ,n8[3]);
    not g224(n516 ,n502);
    nor g225(n245 ,n491 ,n214);
    dff g226(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[5]), .Q(n28[7]));
    not g227(n496 ,n352);
    xor g228(n146 ,n27[2] ,n42[2]);
    not g229(n181 ,n35[1]);
    nor g230(n424 ,n418 ,n422);
    nor g231(n356 ,n188 ,n351);
    or g232(n426 ,n408 ,n423);
    dff g233(.RN(n1), .SN(1'b1), .CK(n0), .D(n158), .Q(n33[1]));
    dff g234(.RN(n1), .SN(1'b1), .CK(n0), .D(n131), .Q(n20[1]));
    dff g235(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[6]), .Q(n24[6]));
    dff g236(.RN(n1), .SN(1'b1), .CK(n0), .D(n57), .Q(n38[0]));
    not g237(n490 ,n16[2]);
    not g238(n54 ,n30[8]);
    not g239(n455 ,n25[3]);
    not g240(n511 ,n1);
    nor g241(n239 ,n181 ,n214);
    xor g242(n177 ,n32[2] ,n167);
    not g243(n481 ,n21[6]);
    not g244(n477 ,n20[0]);
    nor g245(n371 ,n208 ,n367);
    or g246(n328 ,n253 ,n252);
    xor g247(n76 ,n35[0] ,n3[0]);
    or g248(n213 ,n178 ,n205);
    or g249(n61 ,n60 ,n30[13]);
    dff g250(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[0]), .Q(n27[2]));
    xor g251(n96 ,n39[2] ,n9[0]);
    nor g252(n259 ,n432 ,n216);
    dff g253(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[0]), .Q(n26[2]));
    nor g254(n206 ,n37[0] ,n204);
    nor g255(n285 ,n461 ,n215);
    xor g256(n173 ,n118 ,n119);
    dff g257(.RN(n1), .SN(1'b1), .CK(n0), .D(n14[2]), .Q(n14[4]));
    or g258(n400 ,n250 ,n395);
    dff g259(.RN(n1), .SN(1'b1), .CK(n0), .D(n77), .Q(n33[2]));
    not g260(n456 ,n25[6]);
    dff g261(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[5]), .Q(n25[7]));
    xor g262(n134 ,n28[2] ,n40[2]);
    dff g263(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[7]), .Q(n17[7]));
    or g264(n313 ,n277 ,n219);
    not g265(n479 ,n20[1]);
    nor g266(n261 ,n434 ,n209);
    or g267(n305 ,n267 ,n266);
    xnor g268(n112 ,n5[3] ,n36[3]);
    or g269(n309 ,n237 ,n236);
    or g270(n331 ,n303 ,n311);
    nor g271(n282 ,n446 ,n210);
    xor g272(n361 ,n500 ,n36[3]);
    not g273(n520 ,n47[3]);
    dff g274(.RN(n1), .SN(1'b1), .CK(n0), .D(n156), .Q(n25[0]));
    xor g275(n153 ,n26[2] ,n43[2]);
    dff g276(.RN(n1), .SN(1'b1), .CK(n0), .D(n89), .Q(n17[3]));
    or g277(n498 ,n348 ,n346);
    xnor g278(n369 ,n361 ,n35[3]);
    dff g279(.RN(n1), .SN(1'b1), .CK(n0), .D(n141), .Q(n24[2]));
    nor g280(n249 ,n464 ,n212);
    nor g281(n373 ,n208 ,n370);
    dff g282(.RN(n1), .SN(1'b1), .CK(n0), .D(n159), .Q(n33[0]));
    dff g283(.RN(n1), .SN(1'b1), .CK(n0), .D(n162), .Q(n30[2]));
    nor g284(n257 ,n460 ,n216);
    or g285(n321 ,n289 ,n272);
    not g286(n205 ,n204);
    not g287(n517 ,n47[1]);
    xnor g288(n168 ,n74 ,n31[2]);
    nor g289(n365 ,n357 ,n363);
    xor g290(n143 ,n35[1] ,n3[1]);
    not g291(n493 ,n349);
    nor g292(n236 ,n183 ,n212);
    dff g293(.RN(n1), .SN(1'b1), .CK(n0), .D(n14[5]), .Q(n14[7]));
    or g294(n532 ,n527 ,n526);
    xnor g295(n381 ,n376 ,n33[3]);
    nor g296(n357 ,n196 ,n349);
    dff g297(.RN(n1), .SN(1'b1), .CK(n0), .D(n105), .Q(n16[3]));
    xor g298(n104 ,n14[2] ,n46[2]);
    not g299(n468 ,n23[7]);
    or g300(n527 ,n516 ,n515);
    dff g301(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[1]), .Q(n27[3]));
    xnor g302(n114 ,n2[3] ,n3[3]);
    dff g303(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[0]), .Q(n30[8]));
    nor g304(n384 ,n216 ,n381);
    xnor g305(n121 ,n3[3] ,n35[3]);
    xor g306(n80 ,n45[2] ,n7[2]);
    dff g307(.RN(n512), .SN(1'b1), .CK(n0), .D(n507), .Q(n47[1]));
    or g308(n336 ,n302 ,n296);
    xnor g309(n111 ,n2[0] ,n3[0]);
    dff g310(.RN(n512), .SN(1'b1), .CK(n0), .D(n504), .Q(n47[4]));
    not g311(n178 ,n37[0]);
    or g312(n530 ,n522 ,n521);
    or g313(n415 ,n251 ,n409);
    dff g314(.RN(n1), .SN(1'b1), .CK(n0), .D(n84), .Q(n42[3]));
    not g315(n390 ,n389);
    dff g316(.RN(n1), .SN(1'b1), .CK(n0), .D(n137), .Q(n18[3]));
    dff g317(.RN(n1), .SN(1'b1), .CK(n0), .D(n93), .Q(n40[0]));
    dff g318(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[5]), .Q(n26[7]));
    nor g319(n354 ,n208 ,n349);
    nor g320(n276 ,n488 ,n216);
    dff g321(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[4]), .Q(n19[6]));
    xor g322(n171 ,n115 ,n111);
    nor g323(n221 ,n477 ,n208);
    xnor g324(n120 ,n3[2] ,n35[2]);
    xor g325(n150 ,n32[3] ,n31[3]);
    dff g326(.RN(n1), .SN(1'b1), .CK(n0), .D(n496), .Q(n10[7]));
    xnor g327(n119 ,n2[4] ,n3[2]);
    dff g328(.RN(n1), .SN(1'b1), .CK(n0), .D(n38[0]), .Q(n37[0]));
    or g329(n296 ,n257 ,n220);
    not g330(n431 ,n18[1]);
    nor g331(n264 ,n458 ,n215);
    dff g332(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[4]), .Q(n25[6]));
    dff g333(.RN(n1), .SN(1'b1), .CK(n0), .D(n175), .Q(n35[2]));
    xnor g334(n70 ,n8[3] ,n34[3]);
    dff g335(.RN(n1), .SN(1'b1), .CK(n0), .D(n102), .Q(n15[3]));
    xor g336(n100 ,n2[14] ,n3[7]);
    xor g337(n131 ,n19[1] ,n39[1]);
    nor g338(n349 ,n334 ,n339);
    not g339(n188 ,n34[5]);
    not g340(n441 ,n17[6]);
    or g341(n202 ,n179 ,n37[0]);
    dff g342(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[1]), .Q(n30[9]));
    nor g343(n407 ,n209 ,n403);
    xor g344(n101 ,n43[3] ,n4[4]);
    not g345(n57 ,n38[0]);
    xor g346(n151 ,n32[2] ,n31[2]);
    or g347(n521 ,n47[4] ,n47[6]);
    dff g348(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[3]), .Q(n27[5]));
    not g349(n494 ,n351);
    dff g350(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[1]), .Q(n23[3]));
    not g351(n467 ,n22[3]);
    xor g352(n509 ,n38[2] ,n51);
    xnor g353(n158 ,n9[1] ,n69);
    xnor g354(n370 ,n362 ,n35[1]);
    nor g355(n248 ,n492 ,n214);
    dff g356(.RN(n1), .SN(1'b1), .CK(n0), .D(n90), .Q(n34[5]));
    dff g357(.RN(n1), .SN(1'b1), .CK(n0), .D(n91), .Q(n40[2]));
    or g358(n500 ,n345 ,n344);
    dff g359(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[0]), .Q(n25[2]));
    nor g360(n366 ,n356 ,n364);
    or g361(n255 ,n206 ,n207);
    nor g362(n292 ,n185 ,n215);
    or g363(n317 ,n225 ,n280);
    dff g364(.RN(n1), .SN(1'b1), .CK(n0), .D(n85), .Q(n42[2]));
    nor g365(n271 ,n474 ,n215);
    nor g366(n232 ,n470 ,n213);
    not g367(n186 ,n31[2]);
    not g368(n514 ,n508);
    nor g369(n220 ,n484 ,n208);
    nor g370(n281 ,n452 ,n210);
    not g371(n465 ,n23[6]);
    dff g372(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[2]), .Q(n25[4]));
    buf g373(n12[0], 1'b0);
    dff g374(.RN(n1), .SN(1'b1), .CK(n0), .D(n83), .Q(n43[2]));
    not g375(n475 ,n16[7]);
    or g376(n525 ,n517 ,n520);
    nor g377(n237 ,n187 ,n214);
    nor g378(n207 ,n178 ,n199);
    or g379(n533 ,n530 ,n531);
    nor g380(n243 ,n476 ,n214);
    dff g381(.RN(n1), .SN(1'b1), .CK(n0), .D(n14[6]), .Q(n15[6]));
    or g382(n396 ,n372 ,n385);
    nor g383(n241 ,n191 ,n214);
    not g384(n482 ,n22[7]);
    not g385(n449 ,n26[6]);
    xor g386(n87 ,n41[3] ,n6[2]);
    not g387(n194 ,n36[3]);
    dff g388(.RN(n1), .SN(1'b1), .CK(n0), .D(n170), .Q(n35[3]));
    or g389(n338 ,n295 ,n310);
    or g390(n307 ,n270 ,n269);
    or g391(n301 ,n264 ,n263);
    or g392(n394 ,n374 ,n384);
    not g393(n489 ,n17[2]);
    not g394(n478 ,n21[3]);
    dff g395(.RN(n1), .SN(1'b1), .CK(n0), .D(n32[2]), .Q(n11[2]));
    not g396(n458 ,n22[2]);
    nor g397(n267 ,n456 ,n215);
    not g398(n294 ,n293);
    dff g399(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[4]), .Q(n28[6]));
    xor g400(n99 ,n39[0] ,n7[0]);
    dff g401(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[15]), .Q(n14[1]));
    or g402(n406 ,n213 ,n398);
    nor g403(n268 ,n441 ,n210);
    not g404(n483 ,n20[3]);
    dff g405(.RN(n1), .SN(1'b1), .CK(n0), .D(n75), .Q(n33[3]));
    nor g406(n256 ,n481 ,n213);
    nor g407(n226 ,n442 ,n214);
    or g408(n65 ,n53 ,n30[11]);
    xor g409(n135 ,n36[1] ,n5[1]);
    or g410(n364 ,n211 ,n358);
    or g411(n526 ,n513 ,n514);
    dff g412(.RN(n1), .SN(1'b1), .CK(n0), .D(n86), .Q(n42[1]));
    dff g413(.RN(n1), .SN(1'b1), .CK(n0), .D(n498), .Q(n10[1]));
    not g414(n519 ,n47[5]);
    dff g415(.RN(n1), .SN(1'b1), .CK(n0), .D(n98), .Q(n39[1]));
    nor g416(n291 ,n447 ,n216);
    not g417(n435 ,n29[2]);
    nor g418(n385 ,n255 ,n380);
    dff g419(.RN(n1), .SN(1'b1), .CK(n0), .D(n173), .Q(n29[0]));
    not g420(n429 ,n19[7]);
    dff g421(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[3]), .Q(n23[5]));
    nor g422(n409 ,n401 ,n405);
    or g423(n497 ,n341 ,n331);
    nor g424(n289 ,n482 ,n215);
    dff g425(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[1]), .Q(n29[3]));
    dff g426(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[7]), .Q(n30[15]));
    nor g427(n502 ,n37[2] ,n350);
    dff g428(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[7]), .Q(n21[7]));
    dff g429(.RN(n1), .SN(1'b1), .CK(n0), .D(n80), .Q(n45[2]));
    nor g430(n166 ,n66 ,n154);
    xnor g431(n169 ,n70 ,n31[3]);
    not g432(n190 ,n27[3]);
    nor g433(n204 ,n180 ,n37[2]);
    xnor g434(n162 ,n5[2] ,n113);
    dff g435(.RN(n1), .SN(1'b1), .CK(n0), .D(n151), .Q(n31[2]));
    xor g436(n88 ,n41[2] ,n4[2]);
    dff g437(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[7]), .Q(n16[7]));
    nor g438(n273 ,n435 ,n209);
    xnor g439(n164 ,n112 ,n31[3]);
    or g440(n320 ,n246 ,n244);
    dff g441(.RN(n1), .SN(1'b1), .CK(n0), .D(n161), .Q(n30[3]));
    dff g442(.RN(n1), .SN(1'b1), .CK(n0), .D(n78), .Q(n46[2]));
    xor g443(n132 ,n19[0] ,n39[0]);
    xor g444(n84 ,n42[3] ,n6[3]);
    nor g445(n246 ,n439 ,n214);
    dff g446(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[3]), .Q(n25[5]));
    or g447(n152 ,n68 ,n62);
    or g448(n343 ,n316 ,n313);
    dff g449(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[5]), .Q(n19[7]));
    xnor g450(n376 ,n34[3] ,n369);
    nor g451(n355 ,n34[4] ,n493);
    nor g452(n167 ,n63 ,n155);
    not g453(n485 ,n21[7]);
    dff g454(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[4]), .Q(n26[6]));
    not g455(n492 ,n14[7]);
    or g456(n216 ,n178 ,n200);
    or g457(n522 ,n47[0] ,n47[2]);
    or g458(n64 ,n54 ,n30[9]);
    nor g459(n265 ,n466 ,n209);
    nor g460(n228 ,n473 ,n213);
    not g461(n437 ,n18[3]);
    not g462(n443 ,n27[6]);
    not g463(n53 ,n30[12]);
    xnor g464(n411 ,n30[3] ,n404);
    dff g465(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[6]), .Q(n21[6]));
    xor g466(n142 ,n2[7] ,n3[7]);
    not g467(n392 ,n391);
    dff g468(.RN(n1), .SN(1'b1), .CK(n0), .D(n76), .Q(n35[0]));
    or g469(n332 ,n299 ,n297);
    dff g470(.RN(n1), .SN(1'b1), .CK(n0), .D(n145), .Q(n21[1]));
    or g471(n345 ,n320 ,n318);
    xnor g472(n163 ,n5[1] ,n125);
    or g473(n503 ,n353 ,n366);
    or g474(n323 ,n232 ,n286);
    dff g475(.RN(n1), .SN(1'b1), .CK(n0), .D(n101), .Q(n43[3]));
    dff g476(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[2]), .Q(n27[4]));
    dff g477(.RN(n1), .SN(1'b1), .CK(n0), .D(n144), .Q(n24[3]));
    not g478(n515 ,n504);
    nor g479(n227 ,n468 ,n212);
    nor g480(n374 ,n208 ,n369);
    dff g481(.RN(n512), .SN(1'b1), .CK(n0), .D(n503), .Q(n47[5]));
    or g482(n208 ,n37[0] ,n200);
    buf g483(n11[1], 1'b0);
    dff g484(.RN(n1), .SN(1'b1), .CK(n0), .D(n14[7]), .Q(n15[7]));
    dff g485(.RN(n1), .SN(1'b1), .CK(n0), .D(n97), .Q(n23[0]));
    nor g486(n278 ,n436 ,n209);
    nor g487(n258 ,n430 ,n216);
    not g488(n464 ,n23[3]);
    not g489(n187 ,n35[2]);
    not g490(n196 ,n34[4]);
    dff g491(.RN(n1), .SN(1'b1), .CK(n0), .D(n92), .Q(n40[1]));
    nor g492(n238 ,n459 ,n212);
    xor g493(n144 ,n29[3] ,n41[3]);
    dff g494(.RN(n1), .SN(1'b1), .CK(n0), .D(n135), .Q(n36[1]));
    or g495(n427 ,n393 ,n425);
    or g496(n62 ,n56 ,n30[2]);
    or g497(n319 ,n275 ,n223);
    dff g498(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[5]), .Q(n27[7]));
    or g499(n395 ,n373 ,n386);
    not g500(n183 ,n36[2]);
    dff g501(.RN(n1), .SN(1'b1), .CK(n0), .D(n88), .Q(n41[2]));
    not g502(n470 ,n21[1]);
    nor g503(n211 ,n198 ,n204);
    xor g504(n93 ,n40[0] ,n7[1]);
    or g505(n347 ,n324 ,n330);
    nor g506(n287 ,n448 ,n210);
    dff g507(.RN(n1), .SN(1'b1), .CK(n0), .D(n14[4]), .Q(n14[6]));
    dff g508(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[0]), .Q(n19[2]));
    xor g509(n106 ,n23[2] ,n45[2]);
    or g510(n209 ,n37[0] ,n205);
    buf g511(n11[0], 1'b0);
    not g512(n412 ,n411);
    or g513(n302 ,n256 ,n260);
    nor g514(n225 ,n478 ,n213);
    xor g515(n75 ,n33[3] ,n6[3]);
    or g516(n155 ,n64 ,n149);
    nor g517(n402 ,n197 ,n390);
    nor g518(n198 ,n178 ,n37[2]);
    dff g519(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[7]), .Q(n27[1]));
    or g520(n312 ,n245 ,n230);
    nor g521(n351 ,n347 ,n343);
    dff g522(.RN(n1), .SN(1'b1), .CK(n0), .D(n79), .Q(n45[3]));
    or g523(n428 ,n394 ,n426);
    xnor g524(n165 ,n124 ,n31[2]);
    nor g525(n284 ,n467 ,n215);
    not g526(n463 ,n24[6]);
    xnor g527(n382 ,n377 ,n33[1]);
    dff g528(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[1]), .Q(n25[3]));
    xnor g529(n123 ,n2[6] ,n3[3]);
    nor g530(n501 ,n37[2] ,n352);
    xnor g531(n378 ,n34[0] ,n368);
    or g532(n499 ,n333 ,n332);
    or g533(n344 ,n317 ,n314);
    xnor g534(n170 ,n121 ,n32[3]);
    not g535(n195 ,n32[3]);
    xor g536(n91 ,n40[2] ,n9[1]);
    or g537(n425 ,n407 ,n424);
    xnor g538(n377 ,n34[1] ,n370);
    not g539(n512 ,n511);
    or g540(n534 ,n529 ,n532);
    xor g541(n92 ,n40[1] ,n4[1]);
    or g542(n210 ,n37[0] ,n201);
    not g543(n430 ,n28[6]);
    not g544(n59 ,n30[10]);
    or g545(n316 ,n242 ,n278);
    not g546(n48 ,n38[0]);
    nor g547(n218 ,n483 ,n208);
    or g548(n531 ,n528 ,n523);
    nor g549(n386 ,n255 ,n382);
    xor g550(n90 ,n34[5] ,n8[5]);
    nor g551(n417 ,n27[3] ,n411);
    not g552(n433 ,n17[3]);
    dff g553(.RN(n1), .SN(1'b1), .CK(n0), .D(n95), .Q(n39[3]));
    nor g554(n420 ,n190 ,n412);
    nor g555(n423 ,n420 ,n421);
    xnor g556(n388 ,n32[3] ,n381);
    not g557(n473 ,n21[2]);
    or g558(n304 ,n231 ,n265);
    dff g559(.RN(n1), .SN(1'b1), .CK(n0), .D(n100), .Q(n14[0]));
    xor g560(n79 ,n45[3] ,n4[6]);
    not g561(n185 ,n31[3]);
    xor g562(n141 ,n29[2] ,n41[2]);
    not g563(n466 ,n24[7]);
    or g564(n63 ,n59 ,n30[15]);
    xnor g565(n69 ,n6[1] ,n33[1]);
    xnor g566(n117 ,n2[2] ,n3[1]);
    or g567(n342 ,n306 ,n321);
    or g568(n315 ,n274 ,n282);
    or g569(n504 ,n354 ,n365);
    or g570(n67 ,n52 ,n30[4]);
    or g571(n335 ,n309 ,n307);
    dff g572(.RN(n1), .SN(1'b1), .CK(n0), .D(n139), .Q(n24[1]));
    xor g573(n103 ,n34[1] ,n8[1]);
    xnor g574(n116 ,n5[1] ,n8[1]);
    dff g575(.RN(n1), .SN(1'b1), .CK(n0), .D(n509), .Q(n38[2]));
    dff g576(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[1]), .Q(n28[3]));
    dff g577(.RN(n1), .SN(1'b1), .CK(n0), .D(n110), .Q(n41[1]));
    dff g578(.RN(n1), .SN(1'b1), .CK(n0), .D(n494), .Q(n10[5]));
    not g579(n461 ,n25[7]);
    or g580(n507 ,n400 ,n416);
    xor g581(n102 ,n14[3] ,n46[3]);
    or g582(n523 ,n501 ,n507);
    not g583(n189 ,n27[0]);
    dff g584(.RN(n1), .SN(1'b1), .CK(n0), .D(n510), .Q(n38[1]));
    dff g585(.RN(n1), .SN(1'b1), .CK(n0), .D(n150), .Q(n31[3]));
    xor g586(n109 ,n25[2] ,n44[2]);
    dff g587(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[0]), .Q(n28[2]));
    not g588(n476 ,n15[6]);
    or g589(n416 ,n239 ,n410);
    xor g590(n108 ,n25[3] ,n44[3]);
    dff g591(.RN(n1), .SN(1'b1), .CK(n0), .D(n94), .Q(n34[4]));
    not g592(n439 ,n15[3]);
    nor g593(n352 ,n342 ,n337);
    or g594(n297 ,n259 ,n222);
    dff g595(.RN(n512), .SN(1'b1), .CK(n0), .D(n535), .Q(n13));
    dff g596(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[1]), .Q(n19[3]));
    dff g597(.RN(n1), .SN(1'b1), .CK(n0), .D(n106), .Q(n16[2]));
    xnor g598(n413 ,n30[2] ,n403);
    dff g599(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[2]), .Q(n26[4]));
    dff g600(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[6]), .Q(n16[6]));
    xor g601(n172 ,n122 ,n123);
    dff g602(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[4]), .Q(n23[6]));
    not g603(n445 ,n27[7]);
    not g604(n197 ,n27[1]);
    dff g605(.RN(n1), .SN(1'b1), .CK(n0), .D(n104), .Q(n15[2]));
    nor g606(n229 ,n443 ,n213);
    not g607(n49 ,n38[1]);
    xnor g608(n71 ,n6[0] ,n33[0]);
    not g609(n444 ,n16[3]);
    dff g610(.RN(n1), .SN(1'b1), .CK(n0), .D(n497), .Q(n10[0]));
    or g611(n203 ,n178 ,n179);
    dff g612(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[7]), .Q(n20[7]));
    dff g613(.RN(n1), .SN(1'b1), .CK(n0), .D(n138), .Q(n30[5]));
    dff g614(.RN(n1), .SN(1'b1), .CK(n0), .D(n177), .Q(n32[2]));
    not g615(n484 ,n20[6]);
    not g616(n452 ,n26[7]);
    nor g617(n269 ,n182 ,n210);
    nor g618(n235 ,n469 ,n214);
    xnor g619(n125 ,n2[1] ,n3[1]);
    or g620(n300 ,n229 ,n261);
    dff g621(.RN(n1), .SN(1'b1), .CK(n0), .D(n14[0]), .Q(n14[2]));
    dff g622(.RN(n1), .SN(1'b1), .CK(n0), .D(n19[3]), .Q(n19[5]));
    nor g623(n266 ,n449 ,n210);
    dff g624(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[3]), .Q(n26[5]));
    nor g625(n251 ,n184 ,n212);
    dff g626(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[0]), .Q(n29[2]));
    xor g627(n85 ,n42[2] ,n4[3]);
    dff g628(.RN(n1), .SN(1'b1), .CK(n0), .D(n160), .Q(n30[0]));
    nor g629(n263 ,n489 ,n210);
    dff g630(.RN(n1), .SN(1'b1), .CK(n0), .D(n165), .Q(n36[2]));
    dff g631(.RN(n1), .SN(1'b1), .CK(n0), .D(n146), .Q(n21[2]));
    dff g632(.RN(n1), .SN(1'b1), .CK(n0), .D(n32[3]), .Q(n11[3]));
    nor g633(n252 ,n194 ,n212);
    or g634(n311 ,n276 ,n221);
    dff g635(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[4]), .Q(n30[12]));
    dff g636(.RN(n1), .SN(1'b1), .CK(n0), .D(n103), .Q(n34[1]));
    xor g637(n81 ,n44[3] ,n4[5]);
    not g638(n200 ,n199);
    dff g639(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[9]), .Q(n26[1]));
    not g640(n488 ,n18[0]);
    dff g641(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[3]), .Q(n30[11]));
    nor g642(n231 ,n485 ,n213);
    xor g643(n107 ,n34[0] ,n8[0]);
    xor g644(n97 ,n2[12] ,n3[6]);
    nor g645(n358 ,n34[5] ,n494);
    nor g646(n283 ,n433 ,n210);
    xnor g647(n156 ,n8[5] ,n72);
    or g648(n298 ,n258 ,n217);
    not g649(n442 ,n15[7]);
    dff g650(.RN(n1), .SN(1'b1), .CK(n0), .D(n14[1]), .Q(n14[3]));
    nor g651(n244 ,n444 ,n212);
    dff g652(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[1]), .Q(n26[3]));
    or g653(n327 ,n247 ,n249);
    or g654(n337 ,n304 ,n326);
    xor g655(n86 ,n42[1] ,n7[3]);
    not g656(n513 ,n506);
    or g657(n324 ,n248 ,n227);
    xor g658(n129 ,n19[3] ,n39[3]);
    not g659(n191 ,n35[0]);
    nor g660(n250 ,n193 ,n212);
    dff g661(.RN(n1), .SN(1'b1), .CK(n0), .D(n128), .Q(n18[0]));
    dff g662(.RN(n1), .SN(1'b1), .CK(n0), .D(n133), .Q(n30[4]));
    xor g663(n130 ,n19[2] ,n39[2]);
    or g664(n329 ,n235 ,n240);
    dff g665(.RN(n1), .SN(1'b1), .CK(n0), .D(n96), .Q(n39[2]));
    nor g666(n222 ,n480 ,n208);
    not g667(n487 ,n19[6]);
    xor g668(n128 ,n28[0] ,n40[0]);
    dff g669(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[3]), .Q(n29[5]));
    dff g670(.RN(n512), .SN(1'b1), .CK(n0), .D(n502), .Q(n47[6]));
    xnor g671(n389 ,n30[1] ,n382);
    dff g672(.RN(n1), .SN(1'b1), .CK(n0), .D(n147), .Q(n40[3]));
    dff g673(.RN(n1), .SN(1'b1), .CK(n0), .D(n495), .Q(n10[6]));
    dff g674(.RN(n1), .SN(1'b1), .CK(n0), .D(n108), .Q(n22[3]));
    dff g675(.RN(n1), .SN(1'b1), .CK(n0), .D(n132), .Q(n20[0]));
    xor g676(n105 ,n23[3] ,n45[3]);
    xor g677(n138 ,n2[5] ,n3[5]);
    dff g678(.RN(n1), .SN(1'b1), .CK(n0), .D(n99), .Q(n39[0]));
endmodule
