module top(n0, n1, n2, n3);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3;
    wire [7:0] n4;
    wire [7:0] n5;
    wire [3:0] n6;
    wire [15:0] n7;
    wire [15:0] n8;
    wire [31:0] n9;
    wire [63:0] n10;
    wire [7:0] n11;
    wire [3:0] n12;
    wire [7:0] n13;
    wire [3:0] n14;
    wire [15:0] n15;
    wire [3:0] n16;
    wire n17, n18, n19, n20, n21, n22, n23, n24;
    wire n25, n26, n27, n28, n29, n30, n31, n32;
    wire n33, n34, n35, n36, n37, n38, n39, n40;
    wire n41, n42, n43, n44, n45, n46, n47, n48;
    wire n49, n50, n51, n52, n53, n54, n55, n56;
    wire n57, n58, n59, n60, n61, n62, n63, n64;
    wire n65, n66, n67, n68, n69, n70, n71, n72;
    wire n73, n74, n75, n76, n77, n78, n79, n80;
    wire n81, n82, n83, n84, n85, n86, n87, n88;
    wire n89, n90, n91, n92, n93, n94, n95, n96;
    wire n97, n98, n99, n100, n101, n102, n103, n104;
    wire n105, n106, n107, n108, n109, n110, n111, n112;
    wire n113, n114, n115, n116, n117, n118, n119, n120;
    wire n121, n122, n123, n124, n125, n126, n127, n128;
    wire n129, n130, n131, n132, n133, n134, n135, n136;
    wire n137, n138, n139, n140, n141, n142, n143, n144;
    wire n145, n146, n147, n148, n149, n150, n151, n152;
    wire n153, n154, n155, n156, n157, n158, n159, n160;
    wire n161, n162, n163, n164, n165, n166, n167, n168;
    wire n169, n170, n171, n172, n173, n174, n175, n176;
    wire n177, n178, n179, n180, n181, n182, n183, n184;
    wire n185, n186, n187, n188, n189, n190, n191, n192;
    wire n193, n194, n195, n196, n197, n198, n199, n200;
    wire n201, n202, n203, n204, n205, n206, n207, n208;
    wire n209, n210, n211, n212, n213, n214, n215, n216;
    wire n217, n218, n219, n220, n221, n222, n223, n224;
    wire n225, n226, n227, n228, n229, n230, n231, n232;
    wire n233, n234, n235, n236, n237, n238, n239, n240;
    wire n241, n242, n243, n244, n245, n246, n247, n248;
    wire n249, n250, n251, n252, n253, n254, n255, n256;
    wire n257, n258, n259, n260, n261, n262, n263, n264;
    wire n265, n266, n267, n268, n269, n270, n271, n272;
    wire n273, n274, n275, n276, n277, n278, n279, n280;
    wire n281, n282, n283, n284, n285, n286, n287, n288;
    wire n289, n290, n291, n292, n293, n294, n295, n296;
    wire n297, n298, n299, n300, n301, n302, n303, n304;
    wire n305, n306, n307, n308, n309, n310, n311, n312;
    wire n313, n314, n315, n316, n317, n318, n319, n320;
    wire n321, n322, n323, n324, n325, n326, n327, n328;
    wire n329, n330, n331, n332, n333, n334, n335, n336;
    wire n337, n338, n339, n340, n341, n342, n343, n344;
    wire n345, n346, n347, n348, n349, n350, n351, n352;
    wire n353, n354, n355, n356, n357, n358, n359, n360;
    wire n361, n362, n363, n364, n365, n366, n367, n368;
    wire n369, n370, n371, n372, n373, n374, n375, n376;
    wire n377, n378, n379, n380, n381, n382, n383, n384;
    wire n385, n386, n387, n388, n389, n390, n391, n392;
    wire n393, n394, n395, n396, n397, n398, n399, n400;
    wire n401, n402, n403, n404, n405, n406, n407, n408;
    wire n409, n410, n411, n412, n413, n414, n415, n416;
    wire n417, n418, n419, n420, n421, n422, n423, n424;
    wire n425, n426, n427, n428, n429, n430, n431, n432;
    wire n433, n434, n435, n436, n437, n438, n439, n440;
    wire n441, n442, n443, n444, n445, n446, n447, n448;
    wire n449, n450, n451, n452, n453, n454, n455, n456;
    wire n457, n458, n459, n460, n461, n462, n463, n464;
    wire n465, n466, n467, n468, n469, n470, n471, n472;
    wire n473, n474, n475, n476, n477, n478, n479, n480;
    wire n481, n482, n483, n484, n485, n486, n487, n488;
    wire n489, n490, n491, n492, n493, n494, n495, n496;
    wire n497, n498, n499, n500, n501, n502, n503, n504;
    wire n505, n506, n507, n508, n509, n510, n511, n512;
    wire n513, n514, n515, n516, n517, n518, n519, n520;
    wire n521, n522, n523, n524, n525, n526;
    or g0(n322 ,n240 ,n242);
    buf g1(n3[31], n3[63]);
    not g2(n110 ,n109);
    dff g3(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n357), .Q(n8[5]));
    nor g4(n156 ,n133 ,n154);
    not g5(n125 ,n124);
    not g6(n79 ,n15[7]);
    not g7(n225 ,n486);
    nor g8(n265 ,n233 ,n14[0]);
    not g9(n212 ,n496);
    nor g10(n440 ,n236 ,n435);
    not g11(n17 ,n15[6]);
    or g12(n65 ,n58 ,n60);
    nor g13(n422 ,n192 ,n413);
    nor g14(n187 ,n12[1] ,n12[0]);
    not g15(n235 ,n14[0]);
    not g16(n353 ,n354);
    nor g17(n179 ,n8[13] ,n177);
    not g18(n247 ,n15[9]);
    buf g19(n3[32], n3[63]);
    dff g20(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n301), .Q(n5[1]));
    nor g21(n387 ,n192 ,n339);
    nor g22(n365 ,n228 ,n324);
    nor g23(n331 ,n318 ,n271);
    nor g24(n182 ,n8[14] ,n180);
    not g25(n262 ,n15[6]);
    not g26(n263 ,n15[15]);
    nor g27(n438 ,n192 ,n434);
    not g28(n145 ,n144);
    nor g29(n290 ,n233 ,n234);
    not g30(n256 ,n15[2]);
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n381), .Q(n15[6]));
    nor g32(n69 ,n63 ,n67);
    nor g33(n188 ,n184 ,n185);
    not g34(n186 ,n12[2]);
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n391), .Q(n15[13]));
    nor g36(n416 ,n340 ,n388);
    or g37(n25 ,n15[11] ,n15[10]);
    nor g38(n350 ,n234 ,n319);
    nor g39(n519 ,n513 ,n516);
    not g40(n198 ,n488);
    not g41(n116 ,n115);
    not g42(n37 ,n8[3]);
    not g43(n260 ,n15[13]);
    buf g44(n3[0], n3[63]);
    nor g45(n302 ,n255 ,n192);
    nor g46(n418 ,n192 ,n412);
    or g47(n42 ,n8[15] ,n8[14]);
    nor g48(n285 ,n205 ,n462);
    nor g49(n339 ,n312 ,n281);
    nor g50(n520 ,n513 ,n515);
    nor g51(n390 ,n192 ,n344);
    not g52(n254 ,n15[8]);
    or g53(n388 ,n192 ,n354);
    nor g54(n121 ,n86 ,n119);
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n370), .Q(n8[15]));
    not g56(n219 ,n2[2]);
    nor g57(n278 ,n215 ,n462);
    nor g58(n310 ,n257 ,n193);
    not g59(n129 ,n8[13]);
    nor g60(n171 ,n140 ,n169);
    not g61(n85 ,n15[0]);
    buf g62(n3[26], n3[63]);
    not g63(n196 ,n15[14]);
    nor g64(n512 ,n502 ,n510);
    or g65(n267 ,n234 ,n11[0]);
    nor g66(n307 ,n262 ,n193);
    nor g67(n88 ,n80 ,n85);
    or g68(n30 ,n17 ,n28);
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n369), .Q(n8[14]));
    buf g70(n3[44], n3[63]);
    not g71(n251 ,n15[10]);
    nor g72(n312 ,n252 ,n193);
    nor g73(n420 ,n395 ,n409);
    not g74(n101 ,n100);
    nor g75(n340 ,n11[2] ,n290);
    nor g76(n391 ,n192 ,n345);
    not g77(n201 ,n495);
    or g78(n47 ,n40 ,n41);
    or g79(n443 ,n459 ,n4[4]);
    not g80(n236 ,n11[2]);
    nor g81(n467 ,n149 ,n150);
    not g82(n253 ,n15[5]);
    not g83(n77 ,n15[5]);
    xor g84(n437 ,n397 ,n433);
    buf g85(n3[33], n3[63]);
    not g86(n192 ,n1);
    not g87(n514 ,n526);
    buf g88(n3[11], n3[63]);
    nor g89(n432 ,n295 ,n429);
    not g90(n140 ,n8[10]);
    nor g91(n311 ,n256 ,n193);
    nor g92(n165 ,n134 ,n163);
    not g93(n215 ,n498);
    not g94(n460 ,n485);
    nor g95(n105 ,n15[7] ,n103);
    nor g96(n96 ,n15[4] ,n94);
    or g97(n348 ,n464 ,n309);
    or g98(n68 ,n15[15] ,n66);
    nor g99(n103 ,n72 ,n101);
    nor g100(n378 ,n192 ,n330);
    or g101(n453 ,n4[6] ,n452);
    not g102(n137 ,n8[9]);
    xnor g103(n450 ,n447 ,n6[0]);
    xor g104(n481 ,n12[3] ,n191);
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n358), .Q(n8[4]));
    nor g106(n363 ,n460 ,n293);
    nor g107(n346 ,n317 ,n286);
    or g108(n63 ,n56 ,n55);
    not g109(n515 ,n16[2]);
    buf g110(n3[62], n3[63]);
    or g111(n43 ,n8[2] ,n8[0]);
    not g112(n57 ,n15[0]);
    nor g113(n284 ,n207 ,n462);
    nor g114(n375 ,n192 ,n346);
    buf g115(n3[4], n3[63]);
    nor g116(n314 ,n196 ,n193);
    not g117(n74 ,n15[3]);
    or g118(n33 ,n15[7] ,n32);
    nor g119(n176 ,n8[12] ,n174);
    not g120(n104 ,n103);
    or g121(n464 ,n458 ,n456);
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n524), .Q(n16[1]));
    nor g123(n471 ,n161 ,n162);
    nor g124(n487 ,n126 ,n127);
    xor g125(n479 ,n8[15] ,n183);
    nor g126(n300 ,n246 ,n192);
    not g127(n261 ,n4[6]);
    xnor g128(n326 ,n15[0] ,n193);
    buf g129(n3[38], n3[63]);
    buf g130(n3[6], n3[63]);
    not g131(n141 ,n8[0]);
    buf g132(n3[34], n3[63]);
    nor g133(n406 ,n267 ,n348);
    not g134(n216 ,n489);
    buf g135(n3[22], n3[63]);
    nor g136(n127 ,n83 ,n125);
    or g137(n324 ,n192 ,n195);
    nor g138(n337 ,n310 ,n278);
    not g139(n200 ,n500);
    not g140(n222 ,n499);
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n375), .Q(n15[12]));
    buf g142(n3[25], n3[63]);
    buf g143(n3[43], n3[63]);
    xnor g144(n325 ,n526 ,n6[0]);
    not g145(n442 ,n480);
    nor g146(n405 ,n214 ,n353);
    not g147(n429 ,n428);
    buf g148(n3[58], n3[63]);
    nor g149(n100 ,n77 ,n98);
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n523), .Q(n16[2]));
    buf g151(n3[40], n3[63]);
    nor g152(n279 ,n222 ,n462);
    or g153(n264 ,n233 ,n11[1]);
    not g154(n517 ,n16[0]);
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n438), .Q(n10[0]));
    buf g156(n3[50], n3[63]);
    not g157(n203 ,n482);
    nor g158(n270 ,n192 ,n194);
    nor g159(n524 ,n508 ,n509);
    not g160(n18 ,n15[2]);
    or g161(n480 ,n68 ,n71);
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n359), .Q(n8[3]));
    or g163(n441 ,n440 ,n439);
    buf g164(n3[27], n3[63]);
    nor g165(n505 ,n518 ,n2[0]);
    not g166(n231 ,n475);
    nor g167(n120 ,n15[12] ,n118);
    nor g168(n400 ,n240 ,n354);
    nor g169(n347 ,n8[0] ,n324);
    nor g170(n281 ,n200 ,n462);
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n418), .Q(n12[2]));
    not g172(n242 ,n12[3]);
    not g173(n510 ,n509);
    nor g174(n389 ,n192 ,n343);
    not g175(n244 ,n8[0]);
    nor g176(n266 ,n236 ,n11[1]);
    or g177(n415 ,n236 ,n398);
    nor g178(n473 ,n167 ,n168);
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n347), .Q(n8[0]));
    not g180(n113 ,n112);
    nor g181(n272 ,n235 ,n237);
    not g182(n82 ,n15[11]);
    not g183(n189 ,n188);
    nor g184(n411 ,n402 ,n405);
    nor g185(n296 ,n248 ,n192);
    nor g186(n523 ,n511 ,n512);
    nor g187(n292 ,n11[0] ,n11[1]);
    buf g188(n3[3], n3[63]);
    not g189(n195 ,n2[0]);
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n298), .Q(n4[3]));
    not g191(n73 ,n15[13]);
    nor g192(n525 ,n506 ,n505);
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n275), .Q(n4[7]));
    or g194(n427 ,n233 ,n424);
    dff g195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n525), .Q(n16[0]));
    nor g196(n357 ,n208 ,n324);
    not g197(n131 ,n8[4]);
    nor g198(n498 ,n93 ,n94);
    nor g199(n492 ,n111 ,n112);
    buf g200(n3[8], n3[63]);
    not g201(n295 ,n294);
    buf g202(n3[20], n3[63]);
    nor g203(n490 ,n117 ,n118);
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n385), .Q(n15[3]));
    or g205(n349 ,n320 ,n322);
    not g206(n98 ,n97);
    not g207(n259 ,n15[12]);
    or g208(n484 ,n42 ,n53);
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n416), .Q(n14[2]));
    nor g210(n174 ,n138 ,n172);
    or g211(n50 ,n36 ,n49);
    buf g212(n3[42], n3[63]);
    nor g213(n344 ,n314 ,n285);
    buf g214(n3[54], n3[63]);
    not g215(n133 ,n8[5]);
    nor g216(n180 ,n129 ,n178);
    nor g217(n150 ,n130 ,n148);
    nor g218(n271 ,n14[0] ,n463);
    or g219(n70 ,n65 ,n69);
    not g220(n204 ,n479);
    or g221(n320 ,n237 ,n241);
    not g222(n207 ,n492);
    nor g223(n333 ,n306 ,n274);
    xor g224(n455 ,n463 ,n446);
    nor g225(n366 ,n223 ,n324);
    buf g226(n3[51], n3[63]);
    nor g227(n470 ,n158 ,n159);
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n441), .Q(n11[2]));
    not g229(n205 ,n487);
    nor g230(n94 ,n74 ,n92);
    nor g231(n360 ,n221 ,n324);
    nor g232(n408 ,n321 ,n372);
    nor g233(n489 ,n120 ,n121);
    nor g234(n126 ,n15[14] ,n124);
    or g235(n21 ,n15[15] ,n15[14]);
    nor g236(n274 ,n218 ,n462);
    nor g237(n424 ,n220 ,n410);
    nor g238(n287 ,n225 ,n462);
    xor g239(n338 ,n463 ,n7[0]);
    nor g240(n332 ,n305 ,n280);
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n294), .Q(n14[0]));
    buf g242(n3[48], n3[63]);
    nor g243(n273 ,n230 ,n462);
    nor g244(n52 ,n44 ,n51);
    or g245(n58 ,n15[9] ,n15[8]);
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n389), .Q(n15[15]));
    not g247(n239 ,n5[0]);
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n378), .Q(n15[9]));
    nor g249(n93 ,n15[3] ,n91);
    or g250(n23 ,n15[9] ,n15[8]);
    buf g251(n3[52], n3[63]);
    nor g252(n397 ,n192 ,n341);
    not g253(n248 ,n4[4]);
    not g254(n245 ,n15[11]);
    nor g255(n152 ,n8[4] ,n150);
    not g256(n134 ,n8[8]);
    not g257(n246 ,n5[1]);
    xor g258(n3[63] ,n454 ,n455);
    dff g259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n380), .Q(n15[7]));
    or g260(n44 ,n38 ,n39);
    not g261(n502 ,n520);
    dff g262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n366), .Q(n8[10]));
    nor g263(n123 ,n15[13] ,n121);
    not g264(n206 ,n490);
    nor g265(n476 ,n176 ,n177);
    not g266(n220 ,n2[1]);
    not g267(n456 ,n4[3]);
    nor g268(n114 ,n15[10] ,n112);
    dff g269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n361), .Q(n8[1]));
    not g270(n217 ,n470);
    nor g271(n393 ,n462 ,n342);
    not g272(n252 ,n15[1]);
    not g273(n107 ,n106);
    nor g274(n396 ,n192 ,n336);
    nor g275(n495 ,n102 ,n103);
    or g276(n24 ,n15[13] ,n15[12]);
    not g277(n211 ,n465);
    nor g278(n472 ,n164 ,n165);
    nor g279(n359 ,n199 ,n324);
    nor g280(n354 ,n236 ,n291);
    nor g281(n475 ,n173 ,n174);
    or g282(n373 ,n266 ,n350);
    not g283(n221 ,n466);
    nor g284(n430 ,n408 ,n426);
    buf g285(n3[35], n3[63]);
    buf g286(n3[23], n3[63]);
    nor g287(n173 ,n8[11] ,n171);
    not g288(n166 ,n165);
    xor g289(n486 ,n15[15] ,n127);
    not g290(n209 ,n493);
    or g291(n53 ,n47 ,n52);
    not g292(n208 ,n469);
    nor g293(n401 ,n242 ,n354);
    dff g294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n377), .Q(n15[10]));
    nor g295(n28 ,n22 ,n27);
    buf g296(n3[7], n3[63]);
    or g297(n431 ,n192 ,n428);
    or g298(n374 ,n11[2] ,n363);
    nor g299(n351 ,n235 ,n276);
    nor g300(n439 ,n417 ,n436);
    buf g301(n3[19], n3[63]);
    not g302(n154 ,n153);
    nor g303(n328 ,n313 ,n273);
    or g304(n51 ,n45 ,n50);
    buf g305(n3[10], n3[63]);
    not g306(n504 ,n519);
    not g307(n214 ,n483);
    nor g308(n49 ,n8[4] ,n48);
    nor g309(n392 ,n192 ,n353);
    not g310(n78 ,n15[8]);
    not g311(n507 ,n506);
    nor g312(n385 ,n192 ,n337);
    nor g313(n99 ,n15[5] ,n97);
    nor g314(n301 ,n239 ,n192);
    not g315(n240 ,n12[2]);
    nor g316(n468 ,n152 ,n153);
    buf g317(n3[13], n3[63]);
    not g318(n84 ,n15[10]);
    buf g319(n3[16], n3[63]);
    not g320(n202 ,n481);
    nor g321(n404 ,n203 ,n353);
    nor g322(n318 ,n244 ,n235);
    nor g323(n482 ,n190 ,n191);
    nor g324(n377 ,n192 ,n328);
    dff g325(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n270), .Q(n9[0]));
    or g326(n40 ,n8[13] ,n8[12]);
    not g327(n122 ,n121);
    nor g328(n97 ,n75 ,n95);
    dff g329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n390), .Q(n15[14]));
    buf g330(n3[14], n3[63]);
    buf g331(n3[60], n3[63]);
    or g332(n60 ,n15[7] ,n15[6]);
    nor g333(n380 ,n192 ,n333);
    dff g334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n386), .Q(n15[2]));
    nor g335(n518 ,n513 ,n517);
    nor g336(n147 ,n132 ,n145);
    not g337(n157 ,n156);
    dff g338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n365), .Q(n8[9]));
    nor g339(n316 ,n260 ,n193);
    not g340(n291 ,n290);
    not g341(n75 ,n15[4]);
    nor g342(n421 ,n192 ,n411);
    nor g343(n386 ,n192 ,n352);
    nor g344(n323 ,n250 ,n193);
    nor g345(n177 ,n142 ,n175);
    not g346(n19 ,n15[5]);
    dff g347(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n397), .Q(n14[1]));
    nor g348(n399 ,n238 ,n329);
    nor g349(n306 ,n258 ,n193);
    nor g350(n412 ,n400 ,n404);
    or g351(n59 ,n15[13] ,n15[12]);
    buf g352(n3[2], n3[63]);
    or g353(n61 ,n15[11] ,n15[10]);
    not g354(n181 ,n180);
    buf g355(n3[17], n3[63]);
    nor g356(n117 ,n15[11] ,n115);
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n392), .Q(n14[3]));
    not g358(n257 ,n15[3]);
    not g359(n56 ,n15[5]);
    dff g360(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n421), .Q(n12[1]));
    not g361(n238 ,n14[2]);
    nor g362(n112 ,n81 ,n110);
    nor g363(n469 ,n155 ,n156);
    nor g364(n31 ,n19 ,n30);
    not g365(n237 ,n12[0]);
    nor g366(n402 ,n241 ,n354);
    dff g367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n299), .Q(n5[0]));
    nor g368(n368 ,n224 ,n324);
    not g369(n172 ,n171);
    nor g370(n288 ,n206 ,n462);
    xnor g371(n454 ,n451 ,n450);
    not g372(n229 ,n478);
    nor g373(n268 ,n234 ,n480);
    nor g374(n304 ,n247 ,n193);
    not g375(n258 ,n15[7]);
    nor g376(n146 ,n8[2] ,n144);
    nor g377(n521 ,n513 ,n514);
    nor g378(n286 ,n216 ,n462);
    or g379(n410 ,n219 ,n373);
    nor g380(n506 ,n501 ,n503);
    nor g381(n111 ,n15[9] ,n109);
    buf g382(n3[28], n3[63]);
    buf g383(n3[36], n3[63]);
    dff g384(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n379), .Q(n15[8]));
    or g385(n342 ,n11[0] ,n268);
    nor g386(n493 ,n108 ,n109);
    nor g387(n106 ,n79 ,n104);
    nor g388(n282 ,n198 ,n462);
    nor g389(n118 ,n82 ,n116);
    xor g390(n522 ,n521 ,n512);
    not g391(n178 ,n177);
    nor g392(n496 ,n99 ,n100);
    nor g393(n381 ,n192 ,n334);
    dff g394(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n302), .Q(n4[6]));
    xnor g395(n447 ,n7[0] ,n8[0]);
    buf g396(n3[30], n3[63]);
    nor g397(n465 ,n144 ,n143);
    not g398(n516 ,n16[1]);
    not g399(n92 ,n91);
    buf g400(n3[61], n3[63]);
    nor g401(n308 ,n253 ,n193);
    or g402(n22 ,n15[4] ,n15[3]);
    nor g403(n191 ,n186 ,n189);
    or g404(n309 ,n239 ,n243);
    nor g405(n159 ,n128 ,n157);
    nor g406(n413 ,n401 ,n403);
    nor g407(n67 ,n15[2] ,n64);
    nor g408(n474 ,n170 ,n171);
    buf g409(n3[57], n3[63]);
    nor g410(n183 ,n139 ,n181);
    or g411(n409 ,n197 ,n399);
    nor g412(n370 ,n204 ,n324);
    not g413(n76 ,n15[2]);
    nor g414(n153 ,n131 ,n151);
    nor g415(n369 ,n229 ,n324);
    or g416(n276 ,n195 ,n14[2]);
    nor g417(n362 ,n461 ,n291);
    not g418(n55 ,n15[4]);
    nor g419(n275 ,n261 ,n192);
    or g420(n462 ,n443 ,n453);
    not g421(n86 ,n15[12]);
    dff g422(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n300), .Q(n5[2]));
    nor g423(n376 ,n192 ,n327);
    buf g424(n3[41], n3[63]);
    nor g425(n435 ,n432 ,n433);
    or g426(n407 ,n362 ,n374);
    or g427(n341 ,n290 ,n292);
    nor g428(n161 ,n8[7] ,n159);
    not g429(n160 ,n159);
    or g430(n45 ,n35 ,n34);
    not g431(n199 ,n467);
    not g432(n130 ,n8[3]);
    not g433(n503 ,n2[0]);
    buf g434(n3[46], n3[63]);
    nor g435(n508 ,n519 ,n506);
    buf g436(n3[12], n3[63]);
    nor g437(n425 ,n393 ,n415);
    xnor g438(n414 ,n354 ,n12[0]);
    nor g439(n164 ,n8[8] ,n162);
    not g440(n224 ,n477);
    nor g441(n335 ,n308 ,n283);
    not g442(n210 ,n468);
    nor g443(n102 ,n15[6] ,n100);
    not g444(n135 ,n8[7]);
    buf g445(n3[29], n3[63]);
    nor g446(n355 ,n227 ,n324);
    or g447(n26 ,n21 ,n25);
    dff g448(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n384), .Q(n6[0]));
    not g449(n81 ,n15[9]);
    or g450(n463 ,n442 ,n462);
    nor g451(n345 ,n316 ,n282);
    or g452(n29 ,n24 ,n26);
    nor g453(n62 ,n54 ,n57);
    nor g454(n483 ,n188 ,n187);
    not g455(n459 ,n4[5]);
    nor g456(n477 ,n179 ,n180);
    nor g457(n371 ,n231 ,n324);
    not g458(n232 ,n476);
    or g459(n452 ,n5[2] ,n449);
    nor g460(n108 ,n15[8] ,n106);
    buf g461(n3[18], n3[63]);
    not g462(n250 ,n15[4]);
    dff g463(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n269), .Q(n13[0]));
    not g464(n194 ,n526);
    not g465(n233 ,n11[0]);
    dff g466(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n394), .Q(n15[0]));
    not g467(n293 ,n292);
    dff g468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n522), .Q(n526));
    nor g469(n298 ,n243 ,n192);
    nor g470(n299 ,n192 ,n195);
    nor g471(n488 ,n123 ,n124);
    nor g472(n297 ,n249 ,n192);
    nor g473(n398 ,n264 ,n349);
    or g474(n448 ,n5[0] ,n464);
    nor g475(n403 ,n202 ,n353);
    not g476(n80 ,n15[1]);
    nor g477(n90 ,n15[2] ,n88);
    nor g478(n428 ,n425 ,n423);
    not g479(n163 ,n162);
    not g480(n241 ,n12[1]);
    nor g481(n190 ,n12[2] ,n188);
    nor g482(n334 ,n307 ,n289);
    not g483(n136 ,n8[1]);
    not g484(n513 ,n1);
    nor g485(n155 ,n8[5] ,n153);
    or g486(n64 ,n15[3] ,n62);
    nor g487(n367 ,n232 ,n324);
    nor g488(n168 ,n137 ,n166);
    xnor g489(n446 ,n9[0] ,n10[0]);
    buf g490(n3[24], n3[63]);
    dff g491(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n396), .Q(n15[4]));
    or g492(n485 ,n23 ,n33);
    nor g493(n500 ,n88 ,n87);
    not g494(n458 ,n5[1]);
    not g495(n72 ,n15[6]);
    nor g496(n280 ,n209 ,n462);
    nor g497(n343 ,n315 ,n287);
    nor g498(n321 ,n239 ,n238);
    or g499(n71 ,n15[14] ,n70);
    nor g500(n20 ,n15[1] ,n15[0]);
    not g501(n95 ,n94);
    nor g502(n143 ,n8[1] ,n8[0]);
    nor g503(n336 ,n323 ,n277);
    dff g504(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n367), .Q(n8[12]));
    not g505(n255 ,n4[5]);
    nor g506(n315 ,n263 ,n193);
    nor g507(n382 ,n192 ,n335);
    not g508(n175 ,n174);
    not g509(n218 ,n494);
    not g510(n54 ,n15[1]);
    or g511(n32 ,n29 ,n31);
    or g512(n372 ,n14[1] ,n351);
    nor g513(n317 ,n259 ,n193);
    nor g514(n478 ,n182 ,n183);
    nor g515(n303 ,n245 ,n193);
    not g516(n227 ,n471);
    xnor g517(n451 ,n445 ,n444);
    buf g518(n3[5], n3[63]);
    not g519(n38 ,n8[7]);
    nor g520(n379 ,n192 ,n332);
    dff g521(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n376), .Q(n15[11]));
    not g522(n197 ,n14[1]);
    buf g523(n3[49], n3[63]);
    not g524(n249 ,n4[3]);
    nor g525(n423 ,n406 ,n407);
    or g526(n66 ,n59 ,n61);
    nor g527(n361 ,n211 ,n324);
    not g528(n128 ,n8[6]);
    buf g529(n3[39], n3[63]);
    nor g530(n167 ,n8[9] ,n165);
    dff g531(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n371), .Q(n8[11]));
    not g532(n417 ,n416);
    not g533(n193 ,n462);
    buf g534(n3[59], n3[63]);
    nor g535(n494 ,n105 ,n106);
    buf g536(n3[15], n3[63]);
    not g537(n132 ,n8[2]);
    dff g538(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n364), .Q(n8[8]));
    nor g539(n352 ,n311 ,n279);
    not g540(n39 ,n8[6]);
    dff g541(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n356), .Q(n8[6]));
    not g542(n228 ,n473);
    nor g543(n356 ,n217 ,n324);
    not g544(n148 ,n147);
    nor g545(n48 ,n37 ,n46);
    nor g546(n329 ,n272 ,n265);
    not g547(n142 ,n8[12]);
    nor g548(n87 ,n15[1] ,n15[0]);
    nor g549(n124 ,n73 ,n122);
    not g550(n226 ,n497);
    not g551(n184 ,n12[1]);
    nor g552(n294 ,n192 ,n11[0]);
    dff g553(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n422), .Q(n12[3]));
    not g554(n35 ,n8[8]);
    nor g555(n509 ,n504 ,n507);
    buf g556(n3[37], n3[63]);
    nor g557(n395 ,n14[2] ,n331);
    dff g558(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n296), .Q(n4[5]));
    nor g559(n289 ,n201 ,n462);
    not g560(n461 ,n484);
    dff g561(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n297), .Q(n4[4]));
    not g562(n213 ,n472);
    buf g563(n3[9], n3[63]);
    nor g564(n269 ,n235 ,n192);
    buf g565(n3[21], n3[63]);
    nor g566(n358 ,n210 ,n324);
    not g567(n139 ,n8[14]);
    or g568(n41 ,n8[11] ,n8[10]);
    nor g569(n149 ,n8[3] ,n147);
    buf g570(n3[53], n3[63]);
    not g571(n169 ,n168);
    dff g572(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n419), .Q(n12[0]));
    nor g573(n109 ,n78 ,n107);
    dff g574(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n387), .Q(n15[1]));
    not g575(n436 ,n435);
    nor g576(n170 ,n8[10] ,n168);
    not g577(n34 ,n8[5]);
    not g578(n243 ,n5[2]);
    dff g579(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n368), .Q(n8[13]));
    dff g580(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n436), .Q(n11[0]));
    nor g581(n283 ,n212 ,n462);
    nor g582(n277 ,n226 ,n462);
    buf g583(n3[55], n3[63]);
    not g584(n83 ,n15[14]);
    not g585(n223 ,n474);
    dff g586(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n355), .Q(n8[7]));
    nor g587(n499 ,n90 ,n91);
    dff g588(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n382), .Q(n15[5]));
    nor g589(n394 ,n192 ,n326);
    nor g590(n364 ,n213 ,n324);
    nor g591(n491 ,n114 ,n115);
    nor g592(n313 ,n251 ,n193);
    nor g593(n27 ,n18 ,n20);
    not g594(n185 ,n12[0]);
    not g595(n36 ,n8[9]);
    or g596(n426 ,n14[3] ,n420);
    nor g597(n305 ,n254 ,n193);
    nor g598(n115 ,n84 ,n113);
    buf g599(n3[1], n3[63]);
    not g600(n230 ,n491);
    xnor g601(n434 ,n526 ,n430);
    not g602(n119 ,n118);
    not g603(n501 ,n518);
    dff g604(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n360), .Q(n8[2]));
    nor g605(n330 ,n304 ,n284);
    nor g606(n497 ,n96 ,n97);
    buf g607(n3[47], n3[63]);
    nor g608(n384 ,n192 ,n325);
    nor g609(n144 ,n136 ,n141);
    not g610(n457 ,n4[7]);
    nor g611(n162 ,n135 ,n160);
    nor g612(n383 ,n192 ,n338);
    nor g613(n511 ,n520 ,n509);
    nor g614(n466 ,n146 ,n147);
    not g615(n151 ,n150);
    xnor g616(n445 ,n11[0] ,n12[0]);
    buf g617(n3[45], n3[63]);
    nor g618(n419 ,n192 ,n414);
    not g619(n89 ,n88);
    nor g620(n319 ,n236 ,n195);
    nor g621(n91 ,n76 ,n89);
    dff g622(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n383), .Q(n7[0]));
    or g623(n449 ,n457 ,n448);
    nor g624(n327 ,n303 ,n288);
    nor g625(n433 ,n427 ,n431);
    xnor g626(n444 ,n13[0] ,n14[0]);
    dff g627(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n437), .Q(n11[1]));
    nor g628(n46 ,n8[1] ,n43);
    not g629(n138 ,n8[11]);
    not g630(n234 ,n11[1]);
    buf g631(n3[56], n3[63]);
    nor g632(n158 ,n8[6] ,n156);
endmodule
