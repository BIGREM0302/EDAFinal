module top(n0, n1, n7, n8, n9, n2, n3, n4, n5, n14, n15, n6, n16, n17, n10, n11, n12, n13);
    input n0, n1, n2, n3, n4, n5, n6;
    input [6:0] n7;
    input [7:0] n8;
    output [7:0] n9, n10, n11, n12, n13;
    output n14, n15, n16, n17;
    wire n0, n1, n2, n3, n4, n5, n6;
    wire [6:0] n7;
    wire [7:0] n8;
    wire [7:0] n9, n10, n11, n12, n13;
    wire n14, n15, n16, n17;
    wire [2:0] n18;
    wire [4:0] n19;
    wire [4:0] n20;
    wire [3:0] n21;
    wire [15:0] n22;
    wire [7:0] n23;
    wire [7:0] n24;
    wire [7:0] n25;
    wire [7:0] n26;
    wire [7:0] n27;
    wire [7:0] n28;
    wire [7:0] n29;
    wire [7:0] n30;
    wire [7:0] n31;
    wire [7:0] n32;
    wire [7:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [7:0] n36;
    wire [7:0] n37;
    wire [7:0] n38;
    wire [3:0] n39;
    wire [3:0] n40;
    wire [7:0] n41;
    wire [7:0] n42;
    wire [7:0] n43;
    wire [7:0] n44;
    wire [7:0] n45;
    wire [7:0] n46;
    wire [7:0] n47;
    wire [7:0] n48;
    wire [7:0] n49;
    wire [7:0] n50;
    wire [7:0] n51;
    wire [7:0] n52;
    wire [7:0] n53;
    wire [7:0] n54;
    wire [7:0] n55;
    wire [7:0] n56;
    wire [7:0] n57;
    wire [3:0] n58;
    wire [3:0] n59;
    wire [7:0] n60;
    wire n61, n62, n63, n64, n65, n66, n67, n68;
    wire n69, n70, n71, n72, n73, n74, n75, n76;
    wire n77, n78, n79, n80, n81, n82, n83, n84;
    wire n85, n86, n87, n88, n89, n90, n91, n92;
    wire n93, n94, n95, n96, n97, n98, n99, n100;
    wire n101, n102, n103, n104, n105, n106, n107, n108;
    wire n109, n110, n111, n112, n113, n114, n115, n116;
    wire n117, n118, n119, n120, n121, n122, n123, n124;
    wire n125, n126, n127, n128, n129, n130, n131, n132;
    wire n133, n134, n135, n136, n137, n138, n139, n140;
    wire n141, n142, n143, n144, n145, n146, n147, n148;
    wire n149, n150, n151, n152, n153, n154, n155, n156;
    wire n157, n158, n159, n160, n161, n162, n163, n164;
    wire n165, n166, n167, n168, n169, n170, n171, n172;
    wire n173, n174, n175, n176, n177, n178, n179, n180;
    wire n181, n182, n183, n184, n185, n186, n187, n188;
    wire n189, n190, n191, n192, n193, n194, n195, n196;
    wire n197, n198, n199, n200, n201, n202, n203, n204;
    wire n205, n206, n207, n208, n209, n210, n211, n212;
    wire n213, n214, n215, n216, n217, n218, n219, n220;
    wire n221, n222, n223, n224, n225, n226, n227, n228;
    wire n229, n230, n231, n232, n233, n234, n235, n236;
    wire n237, n238, n239, n240, n241, n242, n243, n244;
    wire n245, n246, n247, n248, n249, n250, n251, n252;
    wire n253, n254, n255, n256, n257, n258, n259, n260;
    wire n261, n262, n263, n264, n265, n266, n267, n268;
    wire n269, n270, n271, n272, n273, n274, n275, n276;
    wire n277, n278, n279, n280, n281, n282, n283, n284;
    wire n285, n286, n287, n288, n289, n290, n291, n292;
    wire n293, n294, n295, n296, n297, n298, n299, n300;
    wire n301, n302, n303, n304, n305, n306, n307, n308;
    wire n309, n310, n311, n312, n313, n314, n315, n316;
    wire n317, n318, n319, n320, n321, n322, n323, n324;
    wire n325, n326, n327, n328, n329, n330, n331, n332;
    wire n333, n334, n335, n336, n337, n338, n339, n340;
    wire n341, n342, n343, n344, n345, n346, n347, n348;
    wire n349, n350, n351, n352, n353, n354, n355, n356;
    wire n357, n358, n359, n360, n361, n362, n363, n364;
    wire n365, n366, n367, n368, n369, n370, n371, n372;
    wire n373, n374, n375, n376, n377, n378, n379, n380;
    wire n381, n382, n383, n384, n385, n386, n387, n388;
    wire n389, n390, n391, n392, n393, n394, n395, n396;
    wire n397, n398, n399, n400, n401, n402, n403, n404;
    wire n405, n406, n407, n408, n409, n410, n411, n412;
    wire n413, n414, n415, n416, n417, n418, n419, n420;
    wire n421, n422, n423, n424, n425, n426, n427, n428;
    wire n429, n430, n431, n432, n433, n434, n435, n436;
    wire n437, n438, n439, n440, n441, n442, n443, n444;
    wire n445, n446, n447, n448, n449, n450, n451, n452;
    wire n453, n454, n455, n456, n457, n458, n459, n460;
    wire n461, n462, n463, n464, n465, n466, n467, n468;
    wire n469, n470, n471, n472, n473, n474, n475, n476;
    wire n477, n478, n479, n480, n481, n482, n483, n484;
    wire n485, n486, n487, n488, n489, n490, n491, n492;
    wire n493, n494, n495, n496, n497, n498, n499, n500;
    wire n501, n502, n503, n504, n505, n506, n507, n508;
    wire n509, n510, n511, n512, n513, n514, n515, n516;
    wire n517, n518, n519, n520, n521, n522, n523, n524;
    wire n525, n526, n527, n528, n529, n530, n531, n532;
    wire n533, n534, n535, n536, n537, n538, n539, n540;
    wire n541, n542, n543, n544, n545, n546, n547, n548;
    wire n549, n550, n551, n552, n553, n554, n555, n556;
    wire n557, n558, n559, n560, n561, n562, n563, n564;
    wire n565, n566, n567, n568, n569, n570, n571, n572;
    wire n573, n574, n575, n576, n577, n578, n579, n580;
    wire n581, n582, n583, n584, n585, n586, n587, n588;
    wire n589, n590, n591, n592, n593, n594, n595, n596;
    wire n597, n598, n599, n600, n601, n602, n603, n604;
    wire n605, n606, n607, n608, n609, n610, n611, n612;
    wire n613, n614, n615, n616, n617, n618, n619, n620;
    wire n621, n622, n623, n624, n625, n626, n627, n628;
    wire n629, n630, n631, n632, n633, n634, n635, n636;
    wire n637, n638, n639, n640, n641, n642, n643, n644;
    wire n645, n646, n647, n648, n649, n650, n651, n652;
    wire n653, n654, n655, n656, n657, n658, n659, n660;
    wire n661, n662, n663, n664, n665, n666, n667, n668;
    wire n669, n670, n671, n672, n673, n674, n675, n676;
    wire n677, n678, n679, n680, n681, n682, n683, n684;
    wire n685, n686, n687, n688, n689, n690, n691, n692;
    wire n693, n694, n695, n696, n697, n698, n699, n700;
    wire n701, n702, n703, n704, n705, n706, n707, n708;
    wire n709, n710, n711, n712, n713, n714, n715, n716;
    wire n717, n718, n719, n720, n721, n722, n723, n724;
    wire n725, n726, n727, n728, n729, n730, n731, n732;
    wire n733, n734, n735, n736, n737, n738, n739, n740;
    wire n741, n742, n743, n744, n745, n746, n747, n748;
    wire n749, n750, n751, n752, n753, n754, n755, n756;
    wire n757, n758, n759, n760, n761, n762, n763, n764;
    wire n765, n766, n767, n768, n769, n770, n771, n772;
    wire n773, n774, n775, n776, n777, n778, n779, n780;
    wire n781, n782, n783, n784, n785, n786, n787, n788;
    wire n789, n790, n791, n792, n793, n794, n795, n796;
    wire n797, n798, n799, n800, n801, n802, n803, n804;
    wire n805, n806, n807, n808, n809, n810, n811, n812;
    wire n813, n814, n815, n816, n817, n818, n819, n820;
    wire n821, n822, n823, n824, n825, n826, n827, n828;
    wire n829, n830, n831, n832, n833, n834, n835, n836;
    wire n837, n838, n839, n840, n841, n842, n843, n844;
    wire n845, n846, n847, n848, n849, n850, n851, n852;
    wire n853, n854, n855, n856, n857, n858, n859, n860;
    wire n861, n862, n863, n864, n865, n866, n867, n868;
    wire n869, n870, n871, n872, n873, n874, n875, n876;
    wire n877, n878, n879, n880, n881, n882, n883, n884;
    wire n885, n886, n887, n888, n889, n890, n891, n892;
    wire n893, n894, n895, n896, n897, n898, n899, n900;
    wire n901, n902, n903, n904, n905, n906, n907, n908;
    wire n909, n910, n911, n912, n913, n914, n915, n916;
    wire n917, n918, n919, n920, n921, n922, n923, n924;
    wire n925, n926, n927, n928, n929, n930, n931, n932;
    wire n933, n934, n935, n936, n937, n938, n939, n940;
    wire n941, n942, n943, n944, n945, n946, n947, n948;
    wire n949, n950, n951, n952, n953, n954, n955, n956;
    wire n957, n958, n959, n960, n961, n962, n963, n964;
    wire n965, n966, n967, n968, n969, n970, n971, n972;
    wire n973, n974, n975, n976, n977, n978, n979, n980;
    wire n981, n982, n983, n984, n985, n986, n987, n988;
    wire n989, n990, n991, n992, n993, n994, n995, n996;
    wire n997, n998, n999, n1000, n1001, n1002, n1003, n1004;
    wire n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012;
    wire n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
    wire n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
    wire n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
    wire n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044;
    wire n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052;
    wire n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060;
    wire n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068;
    wire n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076;
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084;
    wire n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092;
    wire n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100;
    wire n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108;
    wire n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116;
    wire n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124;
    wire n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132;
    wire n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140;
    wire n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148;
    wire n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156;
    wire n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164;
    wire n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172;
    wire n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180;
    wire n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188;
    wire n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196;
    wire n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204;
    wire n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
    wire n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220;
    wire n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228;
    wire n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236;
    wire n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244;
    wire n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252;
    wire n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260;
    wire n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268;
    wire n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276;
    wire n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284;
    wire n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292;
    wire n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300;
    wire n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308;
    wire n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;
    wire n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;
    wire n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332;
    wire n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340;
    wire n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348;
    wire n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356;
    wire n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364;
    wire n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372;
    wire n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380;
    wire n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388;
    wire n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396;
    wire n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404;
    wire n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412;
    wire n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420;
    wire n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428;
    wire n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436;
    wire n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444;
    wire n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452;
    wire n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460;
    wire n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468;
    wire n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476;
    wire n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484;
    wire n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492;
    wire n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500;
    wire n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508;
    wire n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516;
    wire n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524;
    wire n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532;
    wire n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540;
    wire n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548;
    wire n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556;
    wire n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564;
    wire n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572;
    wire n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580;
    wire n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588;
    wire n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596;
    wire n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604;
    wire n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612;
    wire n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620;
    wire n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628;
    wire n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636;
    wire n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644;
    wire n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652;
    wire n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660;
    wire n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668;
    wire n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676;
    wire n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684;
    wire n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692;
    wire n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700;
    wire n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708;
    wire n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716;
    wire n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724;
    wire n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732;
    wire n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740;
    wire n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748;
    wire n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756;
    wire n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764;
    wire n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772;
    wire n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780;
    wire n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788;
    wire n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796;
    wire n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804;
    wire n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812;
    wire n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820;
    wire n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828;
    wire n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836;
    wire n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844;
    wire n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852;
    wire n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860;
    wire n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868;
    wire n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876;
    wire n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884;
    wire n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892;
    wire n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900;
    wire n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908;
    wire n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916;
    wire n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924;
    wire n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932;
    wire n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940;
    wire n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948;
    wire n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956;
    wire n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964;
    wire n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972;
    wire n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980;
    wire n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988;
    wire n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996;
    wire n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004;
    wire n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012;
    wire n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020;
    wire n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028;
    wire n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036;
    wire n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044;
    wire n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052;
    wire n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060;
    wire n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068;
    wire n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076;
    wire n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084;
    wire n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092;
    wire n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100;
    wire n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108;
    wire n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116;
    wire n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124;
    wire n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132;
    wire n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140;
    wire n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148;
    wire n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156;
    wire n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164;
    wire n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172;
    wire n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180;
    wire n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188;
    wire n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196;
    wire n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204;
    wire n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212;
    wire n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220;
    wire n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228;
    wire n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236;
    wire n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244;
    wire n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252;
    wire n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260;
    wire n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268;
    wire n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276;
    wire n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284;
    wire n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292;
    wire n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300;
    wire n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308;
    wire n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316;
    wire n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324;
    wire n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332;
    wire n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340;
    wire n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348;
    wire n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356;
    wire n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364;
    wire n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372;
    wire n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380;
    wire n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388;
    wire n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396;
    wire n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404;
    wire n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412;
    wire n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420;
    wire n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428;
    wire n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436;
    wire n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444;
    wire n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452;
    wire n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460;
    wire n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468;
    wire n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476;
    wire n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484;
    wire n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492;
    wire n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500;
    wire n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508;
    wire n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516;
    wire n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524;
    wire n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532;
    wire n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540;
    wire n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548;
    wire n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556;
    wire n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564;
    wire n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572;
    wire n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580;
    wire n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588;
    wire n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596;
    wire n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604;
    wire n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612;
    buf g0(n13[0], n10[0]);
    buf g1(n13[1], n10[1]);
    buf g2(n13[2], n10[0]);
    buf g3(n13[3], n10[1]);
    buf g4(n13[4], n10[6]);
    buf g5(n13[5], n10[7]);
    buf g6(n12[0], n11[0]);
    buf g7(n12[1], n11[1]);
    buf g8(n12[2], n11[2]);
    buf g9(n12[3], 1'b0);
    buf g10(n12[4], 1'b0);
    buf g11(n12[5], 1'b0);
    buf g12(n12[6], 1'b0);
    buf g13(n12[7], 1'b0);
    buf g14(n11[4], 1'b0);
    buf g15(n11[5], 1'b0);
    buf g16(n11[6], 1'b0);
    buf g17(n11[7], 1'b0);
    not g18(n2562 ,n18[0]);
    not g19(n2561 ,n5);
    or g20(n2606 ,n2553 ,n2556);
    or g21(n2605 ,n2555 ,n2560);
    or g22(n2603 ,n2554 ,n2559);
    or g23(n2604 ,n2551 ,n2558);
    or g24(n2602 ,n2552 ,n2557);
    nor g25(n2560 ,n2546 ,n2563);
    nor g26(n2559 ,n2547 ,n2563);
    nor g27(n2558 ,n2542 ,n2563);
    nor g28(n2557 ,n2545 ,n2563);
    nor g29(n2556 ,n2544 ,n2563);
    nor g30(n2555 ,n2540 ,n2550);
    nor g31(n2554 ,n2543 ,n2550);
    nor g32(n2553 ,n2549 ,n2550);
    nor g33(n2552 ,n2548 ,n2550);
    nor g34(n2551 ,n2541 ,n2550);
    not g35(n2563 ,n2550);
    nor g36(n2550 ,n2562 ,n18[1]);
    not g37(n2549 ,n19[4]);
    not g38(n2548 ,n19[0]);
    not g39(n2547 ,n20[1]);
    not g40(n2546 ,n20[3]);
    not g41(n2545 ,n20[0]);
    not g42(n2544 ,n20[4]);
    not g43(n2543 ,n19[1]);
    not g44(n2542 ,n20[2]);
    not g45(n2541 ,n19[2]);
    not g46(n2540 ,n19[3]);
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1641), .Q(n17));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1716), .Q(n21[0]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1713), .Q(n21[1]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1721), .Q(n21[2]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1723), .Q(n21[3]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n700), .Q(n16));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n845), .Q(n22[0]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1559), .Q(n22[1]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1558), .Q(n22[2]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1560), .Q(n22[3]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1561), .Q(n22[4]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1562), .Q(n22[5]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1552), .Q(n22[6]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1543), .Q(n22[7]));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1544), .Q(n22[8]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1545), .Q(n22[9]));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1546), .Q(n22[10]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1547), .Q(n22[11]));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1548), .Q(n22[12]));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1550), .Q(n22[13]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1551), .Q(n22[14]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1549), .Q(n22[15]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n655), .Q(n10[0]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n657), .Q(n10[1]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n654), .Q(n10[6]));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n636), .Q(n10[7]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n622), .Q(n13[6]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n613), .Q(n13[7]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1576), .Q(n11[0]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1575), .Q(n11[1]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n711), .Q(n11[2]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1675), .Q(n11[3]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1938), .Q(n9[0]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1789), .Q(n9[1]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1788), .Q(n9[2]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1787), .Q(n9[3]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1795), .Q(n9[4]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1792), .Q(n9[5]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1794), .Q(n9[6]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1790), .Q(n9[7]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2296), .Q(n23[0]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2217), .Q(n23[1]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2219), .Q(n23[2]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2218), .Q(n23[3]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2216), .Q(n23[4]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2215), .Q(n23[5]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2214), .Q(n23[6]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2213), .Q(n23[7]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2295), .Q(n24[0]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2212), .Q(n24[1]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2211), .Q(n24[2]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2210), .Q(n24[3]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2209), .Q(n24[4]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2208), .Q(n24[5]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2206), .Q(n24[6]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2207), .Q(n24[7]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2406), .Q(n25[0]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2205), .Q(n25[1]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2204), .Q(n25[2]));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2203), .Q(n25[3]));
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2202), .Q(n25[4]));
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2201), .Q(n25[5]));
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2200), .Q(n25[6]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2199), .Q(n25[7]));
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2407), .Q(n26[0]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2198), .Q(n26[1]));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2197), .Q(n26[2]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2196), .Q(n26[3]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2195), .Q(n26[4]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2193), .Q(n26[5]));
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2194), .Q(n26[6]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2192), .Q(n26[7]));
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2408), .Q(n27[0]));
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2191), .Q(n27[1]));
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2190), .Q(n27[2]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2189), .Q(n27[3]));
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2188), .Q(n27[4]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2186), .Q(n27[5]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2185), .Q(n27[6]));
    dff g126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2184), .Q(n27[7]));
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2409), .Q(n28[0]));
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2183), .Q(n28[1]));
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2180), .Q(n28[2]));
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2182), .Q(n28[3]));
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2181), .Q(n28[4]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2179), .Q(n28[5]));
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2178), .Q(n28[6]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2177), .Q(n28[7]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2352), .Q(n29[0]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2176), .Q(n29[1]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2175), .Q(n29[2]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2174), .Q(n29[3]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2173), .Q(n29[4]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2172), .Q(n29[5]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2171), .Q(n29[6]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2170), .Q(n29[7]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2294), .Q(n30[0]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2291), .Q(n30[1]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2293), .Q(n30[2]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2292), .Q(n30[3]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2290), .Q(n30[4]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2289), .Q(n30[5]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2288), .Q(n30[6]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2287), .Q(n30[7]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2309), .Q(n31[0]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2286), .Q(n31[1]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2285), .Q(n31[2]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2284), .Q(n31[3]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2283), .Q(n31[4]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2282), .Q(n31[5]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2281), .Q(n31[6]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2280), .Q(n31[7]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2308), .Q(n32[0]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2279), .Q(n32[1]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2278), .Q(n32[2]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2277), .Q(n32[3]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2276), .Q(n32[4]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2275), .Q(n32[5]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2274), .Q(n32[6]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2273), .Q(n32[7]));
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2307), .Q(n33[0]));
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2271), .Q(n33[1]));
    dff g169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2270), .Q(n33[2]));
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2269), .Q(n33[3]));
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2268), .Q(n33[4]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2267), .Q(n33[5]));
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2265), .Q(n33[6]));
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2266), .Q(n33[7]));
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2306), .Q(n34[0]));
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2264), .Q(n34[1]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2263), .Q(n34[2]));
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2262), .Q(n34[3]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2260), .Q(n34[4]));
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2259), .Q(n34[5]));
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2258), .Q(n34[6]));
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2257), .Q(n34[7]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2305), .Q(n35[0]));
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2256), .Q(n35[1]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2253), .Q(n35[2]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2251), .Q(n35[3]));
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2246), .Q(n35[4]));
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2250), .Q(n35[5]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2248), .Q(n35[6]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2187), .Q(n35[7]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2304), .Q(n36[0]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2245), .Q(n36[1]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2244), .Q(n36[2]));
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2242), .Q(n36[3]));
    dff g195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2241), .Q(n36[4]));
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2240), .Q(n36[5]));
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2238), .Q(n36[6]));
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2252), .Q(n36[7]));
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2303), .Q(n37[0]));
    dff g200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2272), .Q(n37[1]));
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2236), .Q(n37[2]));
    dff g202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2229), .Q(n37[3]));
    dff g203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2234), .Q(n37[4]));
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2233), .Q(n37[5]));
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2232), .Q(n37[6]));
    dff g206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2231), .Q(n37[7]));
    dff g207(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2302), .Q(n38[0]));
    dff g208(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2249), .Q(n38[1]));
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2230), .Q(n38[2]));
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2228), .Q(n38[3]));
    dff g211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2226), .Q(n38[4]));
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2239), .Q(n38[5]));
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2225), .Q(n38[6]));
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2224), .Q(n38[7]));
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2223), .Q(n20[0]));
    dff g216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2301), .Q(n20[1]));
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2300), .Q(n20[2]));
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2299), .Q(n20[3]));
    dff g219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2298), .Q(n20[4]));
    dff g220(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n756), .Q(n39[0]));
    dff g221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1427), .Q(n39[1]));
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1426), .Q(n39[2]));
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1425), .Q(n39[3]));
    dff g224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1717), .Q(n40[0]));
    dff g225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2220), .Q(n40[1]));
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2222), .Q(n40[2]));
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2221), .Q(n40[3]));
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1640), .Q(n41[0]));
    dff g229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1633), .Q(n41[1]));
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1632), .Q(n41[2]));
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1631), .Q(n41[3]));
    dff g232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1630), .Q(n41[4]));
    dff g233(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1629), .Q(n41[5]));
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1628), .Q(n41[6]));
    dff g235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1627), .Q(n41[7]));
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1639), .Q(n14));
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2417), .Q(n15));
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1784), .Q(n18[0]));
    dff g239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1980), .Q(n18[1]));
    dff g240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1786), .Q(n18[2]));
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n706), .Q(n10[2]));
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n707), .Q(n10[3]));
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n701), .Q(n10[4]));
    dff g244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n702), .Q(n10[5]));
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1454), .Q(n42[0]));
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1419), .Q(n42[1]));
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1418), .Q(n42[2]));
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1417), .Q(n42[3]));
    dff g249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1416), .Q(n42[4]));
    dff g250(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1415), .Q(n42[5]));
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1414), .Q(n42[6]));
    dff g252(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1413), .Q(n42[7]));
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1453), .Q(n43[0]));
    dff g254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1412), .Q(n43[1]));
    dff g255(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1411), .Q(n43[2]));
    dff g256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1410), .Q(n43[3]));
    dff g257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1409), .Q(n43[4]));
    dff g258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1408), .Q(n43[5]));
    dff g259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1406), .Q(n43[6]));
    dff g260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1405), .Q(n43[7]));
    dff g261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1452), .Q(n44[0]));
    dff g262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1404), .Q(n44[1]));
    dff g263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1403), .Q(n44[2]));
    dff g264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1402), .Q(n44[3]));
    dff g265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1401), .Q(n44[4]));
    dff g266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1400), .Q(n44[5]));
    dff g267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1398), .Q(n44[6]));
    dff g268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1397), .Q(n44[7]));
    dff g269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1451), .Q(n45[0]));
    dff g270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1396), .Q(n45[1]));
    dff g271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1395), .Q(n45[2]));
    dff g272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1394), .Q(n45[3]));
    dff g273(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1393), .Q(n45[4]));
    dff g274(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1392), .Q(n45[5]));
    dff g275(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1391), .Q(n45[6]));
    dff g276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1390), .Q(n45[7]));
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1450), .Q(n46[0]));
    dff g278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1435), .Q(n46[1]));
    dff g279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1388), .Q(n46[2]));
    dff g280(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1387), .Q(n46[3]));
    dff g281(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1386), .Q(n46[4]));
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1385), .Q(n46[5]));
    dff g283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1384), .Q(n46[6]));
    dff g284(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1383), .Q(n46[7]));
    dff g285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1449), .Q(n47[0]));
    dff g286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1382), .Q(n47[1]));
    dff g287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1381), .Q(n47[2]));
    dff g288(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1380), .Q(n47[3]));
    dff g289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1379), .Q(n47[4]));
    dff g290(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1378), .Q(n47[5]));
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1377), .Q(n47[6]));
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1376), .Q(n47[7]));
    dff g293(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1448), .Q(n48[0]));
    dff g294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1375), .Q(n48[1]));
    dff g295(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1374), .Q(n48[2]));
    dff g296(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1373), .Q(n48[3]));
    dff g297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1372), .Q(n48[4]));
    dff g298(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1432), .Q(n48[5]));
    dff g299(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1371), .Q(n48[6]));
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1370), .Q(n48[7]));
    dff g301(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1446), .Q(n49[0]));
    dff g302(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1369), .Q(n49[1]));
    dff g303(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1368), .Q(n49[2]));
    dff g304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1367), .Q(n49[3]));
    dff g305(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1366), .Q(n49[4]));
    dff g306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1365), .Q(n49[5]));
    dff g307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1364), .Q(n49[6]));
    dff g308(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1363), .Q(n49[7]));
    dff g309(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1457), .Q(n50[0]));
    dff g310(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1362), .Q(n50[1]));
    dff g311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1361), .Q(n50[2]));
    dff g312(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1360), .Q(n50[3]));
    dff g313(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1359), .Q(n50[4]));
    dff g314(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1358), .Q(n50[5]));
    dff g315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1357), .Q(n50[6]));
    dff g316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1356), .Q(n50[7]));
    dff g317(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1445), .Q(n51[0]));
    dff g318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1353), .Q(n51[1]));
    dff g319(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1433), .Q(n51[2]));
    dff g320(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1352), .Q(n51[3]));
    dff g321(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1349), .Q(n51[4]));
    dff g322(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1354), .Q(n51[5]));
    dff g323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1351), .Q(n51[6]));
    dff g324(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1350), .Q(n51[7]));
    dff g325(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1447), .Q(n52[0]));
    dff g326(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1348), .Q(n52[1]));
    dff g327(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1347), .Q(n52[2]));
    dff g328(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1399), .Q(n52[3]));
    dff g329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1346), .Q(n52[4]));
    dff g330(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1345), .Q(n52[5]));
    dff g331(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1423), .Q(n52[6]));
    dff g332(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1428), .Q(n52[7]));
    dff g333(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1444), .Q(n53[0]));
    dff g334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1443), .Q(n53[1]));
    dff g335(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1431), .Q(n53[2]));
    dff g336(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1442), .Q(n53[3]));
    dff g337(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1441), .Q(n53[4]));
    dff g338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1440), .Q(n53[5]));
    dff g339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1439), .Q(n53[6]));
    dff g340(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1438), .Q(n53[7]));
    dff g341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1460), .Q(n54[0]));
    dff g342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1455), .Q(n54[1]));
    dff g343(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1434), .Q(n54[2]));
    dff g344(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1469), .Q(n54[3]));
    dff g345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1476), .Q(n54[4]));
    dff g346(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1478), .Q(n54[5]));
    dff g347(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1462), .Q(n54[6]));
    dff g348(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1491), .Q(n54[7]));
    dff g349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1456), .Q(n55[0]));
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1502), .Q(n55[1]));
    dff g351(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1508), .Q(n55[2]));
    dff g352(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1509), .Q(n55[3]));
    dff g353(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1355), .Q(n55[4]));
    dff g354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1510), .Q(n55[5]));
    dff g355(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1511), .Q(n55[6]));
    dff g356(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1420), .Q(n55[7]));
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1458), .Q(n56[0]));
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1512), .Q(n56[1]));
    dff g359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1407), .Q(n56[2]));
    dff g360(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1513), .Q(n56[3]));
    dff g361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1514), .Q(n56[4]));
    dff g362(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1429), .Q(n56[5]));
    dff g363(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1430), .Q(n56[6]));
    dff g364(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1389), .Q(n56[7]));
    dff g365(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1210), .Q(n57[0]));
    dff g366(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1173), .Q(n57[1]));
    dff g367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1184), .Q(n57[2]));
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1178), .Q(n57[3]));
    dff g369(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1183), .Q(n57[4]));
    dff g370(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1164), .Q(n57[5]));
    dff g371(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1182), .Q(n57[6]));
    dff g372(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1188), .Q(n57[7]));
    dff g373(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2064), .Q(n19[0]));
    dff g374(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1984), .Q(n19[1]));
    dff g375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1983), .Q(n19[2]));
    dff g376(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1982), .Q(n19[3]));
    dff g377(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1981), .Q(n19[4]));
    dff g378(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1783), .Q(n58[0]));
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1975), .Q(n58[1]));
    dff g380(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1974), .Q(n58[2]));
    dff g381(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1973), .Q(n58[3]));
    dff g382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n786), .Q(n59[0]));
    dff g383(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n843), .Q(n59[1]));
    dff g384(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n841), .Q(n59[2]));
    dff g385(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n842), .Q(n59[3]));
    dff g386(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2530), .Q(n60[0]));
    dff g387(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2539), .Q(n60[1]));
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2534), .Q(n60[2]));
    dff g389(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2538), .Q(n60[3]));
    dff g390(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2537), .Q(n60[4]));
    dff g391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2535), .Q(n60[5]));
    dff g392(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2536), .Q(n60[6]));
    dff g393(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2533), .Q(n60[7]));
    or g394(n2539 ,n1953 ,n2532);
    or g395(n2538 ,n1949 ,n2529);
    or g396(n2537 ,n1943 ,n2526);
    or g397(n2536 ,n1945 ,n2528);
    or g398(n2535 ,n1946 ,n2527);
    or g399(n2534 ,n1951 ,n2531);
    or g400(n2533 ,n1942 ,n2525);
    or g401(n2532 ,n1611 ,n2523);
    or g402(n2531 ,n1614 ,n2524);
    or g403(n2530 ,n2416 ,n2522);
    or g404(n2529 ,n1609 ,n2521);
    or g405(n2528 ,n1610 ,n2520);
    or g406(n2527 ,n1612 ,n2519);
    or g407(n2526 ,n1622 ,n2518);
    or g408(n2525 ,n1608 ,n2517);
    or g409(n2524 ,n2379 ,n2516);
    or g410(n2523 ,n2390 ,n2515);
    or g411(n2522 ,n201 ,n2514);
    or g412(n2521 ,n2367 ,n2513);
    or g413(n2520 ,n2330 ,n2512);
    or g414(n2519 ,n2342 ,n2511);
    or g415(n2518 ,n2354 ,n2510);
    or g416(n2517 ,n2320 ,n2509);
    or g417(n2516 ,n2477 ,n2508);
    or g418(n2515 ,n2480 ,n2507);
    or g419(n2514 ,n2483 ,n2506);
    or g420(n2513 ,n2474 ,n2505);
    or g421(n2512 ,n2466 ,n2504);
    or g422(n2511 ,n2469 ,n2503);
    or g423(n2510 ,n2472 ,n2502);
    or g424(n2509 ,n2463 ,n2501);
    or g425(n2508 ,n2427 ,n2500);
    or g426(n2507 ,n2420 ,n2499);
    or g427(n2506 ,n2414 ,n2498);
    or g428(n2505 ,n2433 ,n2497);
    or g429(n2504 ,n2451 ,n2496);
    or g430(n2503 ,n2445 ,n2495);
    or g431(n2502 ,n2439 ,n2494);
    or g432(n2501 ,n2457 ,n2493);
    or g433(n2500 ,n2375 ,n2492);
    or g434(n2499 ,n2386 ,n2491);
    or g435(n2498 ,n2400 ,n2490);
    or g436(n2497 ,n2363 ,n2489);
    or g437(n2496 ,n2326 ,n2488);
    or g438(n2495 ,n2338 ,n2487);
    or g439(n2494 ,n2350 ,n2486);
    or g440(n2493 ,n2317 ,n2485);
    or g441(n2492 ,n2476 ,n2475);
    or g442(n2491 ,n2479 ,n2484);
    or g443(n2490 ,n2482 ,n2481);
    or g444(n2489 ,n2478 ,n2473);
    or g445(n2488 ,n2465 ,n2464);
    or g446(n2487 ,n2468 ,n2467);
    or g447(n2486 ,n2471 ,n2470);
    or g448(n2485 ,n2462 ,n2461);
    or g449(n2484 ,n2423 ,n2424);
    or g450(n2483 ,n2415 ,n2261);
    or g451(n2482 ,n2413 ,n2412);
    or g452(n2481 ,n2411 ,n2418);
    or g453(n2480 ,n2419 ,n2255);
    or g454(n2479 ,n2421 ,n2422);
    or g455(n2478 ,n2434 ,n2435);
    or g456(n2477 ,n2426 ,n2247);
    or g457(n2476 ,n2428 ,n2429);
    or g458(n2475 ,n2430 ,n2431);
    or g459(n2474 ,n2432 ,n2243);
    or g460(n2473 ,n2436 ,n2437);
    or g461(n2472 ,n2438 ,n2237);
    or g462(n2471 ,n2440 ,n2441);
    or g463(n2470 ,n2443 ,n2442);
    or g464(n2469 ,n2444 ,n2235);
    or g465(n2468 ,n2446 ,n2447);
    or g466(n2467 ,n2448 ,n2449);
    or g467(n2466 ,n2450 ,n2254);
    or g468(n2465 ,n2452 ,n2453);
    or g469(n2464 ,n2454 ,n2455);
    or g470(n2463 ,n2456 ,n2227);
    or g471(n2462 ,n2425 ,n2458);
    or g472(n2461 ,n2459 ,n2460);
    or g473(n2460 ,n2312 ,n2355);
    or g474(n2459 ,n2087 ,n2313);
    or g475(n2458 ,n2368 ,n2314);
    or g476(n2457 ,n2318 ,n2391);
    or g477(n2456 ,n2077 ,n2319);
    or g478(n2455 ,n2321 ,n2377);
    or g479(n2454 ,n2114 ,n2322);
    or g480(n2453 ,n2346 ,n2323);
    or g481(n2452 ,n2324 ,n2325);
    or g482(n2451 ,n2328 ,n2327);
    or g483(n2450 ,n2169 ,n2329);
    or g484(n2449 ,n2332 ,n2331);
    or g485(n2448 ,n2153 ,n2333);
    or g486(n2447 ,n2336 ,n2335);
    or g487(n2446 ,n2337 ,n2334);
    or g488(n2445 ,n2340 ,n2339);
    or g489(n2444 ,n2084 ,n2341);
    or g490(n2443 ,n2088 ,n2345);
    or g491(n2442 ,n2343 ,n2344);
    or g492(n2441 ,n2347 ,n2405);
    or g493(n2440 ,n2349 ,n2348);
    or g494(n2439 ,n2410 ,n2351);
    or g495(n2438 ,n2092 ,n2353);
    or g496(n2437 ,n2357 ,n2356);
    or g497(n2436 ,n2061 ,n2358);
    or g498(n2435 ,n2360 ,n2359);
    or g499(n2434 ,n2362 ,n2361);
    or g500(n2433 ,n2365 ,n2364);
    or g501(n2432 ,n2099 ,n2366);
    or g502(n2431 ,n2369 ,n2311);
    or g503(n2430 ,n2033 ,n2370);
    or g504(n2429 ,n2373 ,n2372);
    or g505(n2428 ,n2371 ,n2374);
    or g506(n2427 ,n2376 ,n2310);
    or g507(n2426 ,n2105 ,n2378);
    or g508(n2425 ,n2315 ,n2316);
    or g509(n2424 ,n2381 ,n2380);
    or g510(n2423 ,n2109 ,n2382);
    or g511(n2422 ,n2383 ,n2393);
    or g512(n2421 ,n2385 ,n2384);
    or g513(n2420 ,n2387 ,n2388);
    or g514(n2419 ,n2112 ,n2389);
    or g515(n2418 ,n2394 ,n2392);
    or g516(n2417 ,n1231 ,n2297);
    or g517(n2416 ,n1955 ,n2404);
    or g518(n2415 ,n2123 ,n2403);
    or g519(n2414 ,n2402 ,n2401);
    or g520(n2413 ,n2399 ,n2398);
    or g521(n2412 ,n2397 ,n2396);
    or g522(n2411 ,n2116 ,n2395);
    nor g523(n2410 ,n442 ,n2068);
    or g524(n2409 ,n2015 ,n1995);
    or g525(n2408 ,n2024 ,n1994);
    or g526(n2407 ,n2032 ,n1993);
    or g527(n2406 ,n2041 ,n1992);
    nor g528(n2405 ,n318 ,n2073);
    nor g529(n2404 ,n498 ,n2065);
    nor g530(n2403 ,n487 ,n2067);
    nor g531(n2402 ,n467 ,n2068);
    nor g532(n2401 ,n271 ,n2069);
    nor g533(n2400 ,n236 ,n2076);
    nor g534(n2399 ,n337 ,n2066);
    nor g535(n2398 ,n511 ,n2071);
    nor g536(n2397 ,n547 ,n2072);
    nor g537(n2396 ,n576 ,n2073);
    nor g538(n2395 ,n485 ,n2075);
    nor g539(n2394 ,n239 ,n2070);
    nor g540(n2393 ,n534 ,n2073);
    nor g541(n2392 ,n549 ,n2074);
    nor g542(n2391 ,n577 ,n2069);
    nor g543(n2390 ,n447 ,n2065);
    nor g544(n2389 ,n310 ,n2067);
    nor g545(n2388 ,n473 ,n2069);
    nor g546(n2387 ,n254 ,n2068);
    nor g547(n2386 ,n272 ,n2076);
    nor g548(n2385 ,n595 ,n2066);
    nor g549(n2384 ,n452 ,n2071);
    nor g550(n2383 ,n535 ,n2072);
    nor g551(n2382 ,n565 ,n2075);
    nor g552(n2381 ,n491 ,n2070);
    nor g553(n2380 ,n268 ,n2074);
    nor g554(n2379 ,n322 ,n2065);
    nor g555(n2378 ,n540 ,n2067);
    nor g556(n2377 ,n568 ,n2074);
    nor g557(n2376 ,n465 ,n2068);
    nor g558(n2375 ,n554 ,n2076);
    nor g559(n2374 ,n346 ,n2071);
    nor g560(n2373 ,n569 ,n2072);
    nor g561(n2372 ,n470 ,n2073);
    nor g562(n2371 ,n482 ,n2066);
    nor g563(n2370 ,n538 ,n2075);
    nor g564(n2369 ,n599 ,n2070);
    nor g565(n2368 ,n471 ,n2072);
    nor g566(n2367 ,n326 ,n2065);
    nor g567(n2366 ,n286 ,n2067);
    nor g568(n2365 ,n523 ,n2068);
    nor g569(n2364 ,n446 ,n2069);
    nor g570(n2363 ,n558 ,n2076);
    nor g571(n2362 ,n323 ,n2066);
    nor g572(n2361 ,n469 ,n2071);
    nor g573(n2360 ,n308 ,n2072);
    nor g574(n2359 ,n460 ,n2073);
    nor g575(n2358 ,n288 ,n2075);
    nor g576(n2357 ,n453 ,n2070);
    nor g577(n2356 ,n548 ,n2074);
    nor g578(n2355 ,n496 ,n2074);
    nor g579(n2354 ,n591 ,n2065);
    nor g580(n2353 ,n325 ,n2067);
    or g581(n2352 ,n2007 ,n1996);
    nor g582(n2351 ,n594 ,n2069);
    nor g583(n2350 ,n528 ,n2076);
    nor g584(n2349 ,n531 ,n2066);
    nor g585(n2348 ,n529 ,n2071);
    nor g586(n2347 ,n483 ,n2072);
    nor g587(n2346 ,n501 ,n2072);
    nor g588(n2345 ,n502 ,n2075);
    nor g589(n2344 ,n600 ,n2074);
    nor g590(n2343 ,n303 ,n2070);
    nor g591(n2342 ,n457 ,n2065);
    nor g592(n2341 ,n354 ,n2067);
    nor g593(n2340 ,n449 ,n2068);
    nor g594(n2339 ,n592 ,n2069);
    nor g595(n2338 ,n537 ,n2076);
    nor g596(n2337 ,n484 ,n2066);
    nor g597(n2336 ,n295 ,n2072);
    nor g598(n2335 ,n266 ,n2073);
    nor g599(n2334 ,n557 ,n2071);
    nor g600(n2333 ,n258 ,n2075);
    nor g601(n2332 ,n315 ,n2070);
    nor g602(n2331 ,n597 ,n2074);
    nor g603(n2330 ,n311 ,n2065);
    nor g604(n2329 ,n486 ,n2067);
    nor g605(n2328 ,n532 ,n2068);
    nor g606(n2327 ,n536 ,n2069);
    nor g607(n2326 ,n476 ,n2076);
    nor g608(n2325 ,n445 ,n2071);
    nor g609(n2324 ,n468 ,n2066);
    nor g610(n2323 ,n277 ,n2073);
    nor g611(n2322 ,n455 ,n2075);
    nor g612(n2321 ,n459 ,n2070);
    nor g613(n2320 ,n334 ,n2065);
    nor g614(n2319 ,n480 ,n2067);
    nor g615(n2318 ,n290 ,n2068);
    nor g616(n2317 ,n296 ,n2076);
    nor g617(n2316 ,n593 ,n2071);
    nor g618(n2315 ,n248 ,n2066);
    nor g619(n2314 ,n280 ,n2073);
    nor g620(n2313 ,n596 ,n2075);
    nor g621(n2312 ,n514 ,n2070);
    nor g622(n2311 ,n464 ,n2074);
    nor g623(n2310 ,n500 ,n2069);
    or g624(n2309 ,n2151 ,n1978);
    or g625(n2308 ,n2143 ,n1977);
    or g626(n2307 ,n2133 ,n1976);
    or g627(n2306 ,n2125 ,n1972);
    or g628(n2305 ,n2113 ,n1987);
    or g629(n2304 ,n2101 ,n1986);
    or g630(n2303 ,n2115 ,n1988);
    or g631(n2302 ,n2168 ,n1989);
    or g632(n2301 ,n2162 ,n1671);
    or g633(n2300 ,n2161 ,n1673);
    or g634(n2299 ,n2160 ,n1677);
    or g635(n2298 ,n1998 ,n1678);
    or g636(n2297 ,n1685 ,n1985);
    or g637(n2296 ,n2058 ,n1990);
    or g638(n2295 ,n2049 ,n1991);
    or g639(n2294 ,n1999 ,n1979);
    or g640(n2293 ,n1914 ,n2158);
    or g641(n2292 ,n1913 ,n2157);
    or g642(n2291 ,n1915 ,n2159);
    or g643(n2290 ,n1912 ,n2156);
    or g644(n2289 ,n1911 ,n2155);
    or g645(n2288 ,n1909 ,n2154);
    or g646(n2287 ,n1932 ,n2152);
    or g647(n2286 ,n1907 ,n2150);
    or g648(n2285 ,n1906 ,n2149);
    or g649(n2284 ,n1905 ,n2148);
    or g650(n2283 ,n1904 ,n2147);
    or g651(n2282 ,n1903 ,n2146);
    or g652(n2281 ,n1902 ,n2145);
    or g653(n2280 ,n1931 ,n2144);
    or g654(n2279 ,n1900 ,n2141);
    or g655(n2278 ,n1899 ,n2140);
    or g656(n2277 ,n1898 ,n2138);
    or g657(n2276 ,n1897 ,n2137);
    or g658(n2275 ,n1896 ,n2136);
    or g659(n2274 ,n1895 ,n2135);
    or g660(n2273 ,n1930 ,n2134);
    or g661(n2272 ,n1892 ,n2086);
    or g662(n2271 ,n1893 ,n2132);
    or g663(n2270 ,n1889 ,n2131);
    or g664(n2269 ,n1791 ,n2130);
    or g665(n2268 ,n1891 ,n2129);
    or g666(n2267 ,n1880 ,n2127);
    or g667(n2266 ,n1929 ,n2126);
    or g668(n2265 ,n1963 ,n2128);
    or g669(n2264 ,n1887 ,n2124);
    or g670(n2263 ,n1881 ,n2122);
    or g671(n2262 ,n1886 ,n2120);
    or g672(n2261 ,n2121 ,n1954);
    or g673(n2260 ,n1885 ,n2119);
    or g674(n2259 ,n1883 ,n2118);
    or g675(n2258 ,n1882 ,n2117);
    or g676(n2257 ,n1925 ,n2079);
    or g677(n2256 ,n1939 ,n2111);
    or g678(n2255 ,n2096 ,n1952);
    or g679(n2254 ,n2167 ,n1944);
    or g680(n2253 ,n1935 ,n2110);
    or g681(n2252 ,n1927 ,n2089);
    or g682(n2251 ,n1941 ,n2107);
    or g683(n2250 ,n1878 ,n2103);
    or g684(n2249 ,n1801 ,n1997);
    or g685(n2248 ,n1818 ,n2016);
    or g686(n2247 ,n2104 ,n1950);
    or g687(n2246 ,n1804 ,n2106);
    or g688(n2245 ,n1844 ,n2100);
    or g689(n2244 ,n1855 ,n2098);
    or g690(n2243 ,n2051 ,n1948);
    or g691(n2242 ,n1936 ,n2081);
    or g692(n2241 ,n1966 ,n2095);
    or g693(n2240 ,n1890 ,n2093);
    or g694(n2239 ,n1799 ,n2062);
    or g695(n2238 ,n1856 ,n2091);
    or g696(n2237 ,n2090 ,n1947);
    or g697(n2236 ,n1962 ,n2085);
    or g698(n2235 ,n2139 ,n1957);
    or g699(n2234 ,n1964 ,n2082);
    or g700(n2233 ,n1879 ,n2080);
    or g701(n2232 ,n1884 ,n2078);
    or g702(n2231 ,n1926 ,n2097);
    or g703(n2230 ,n1800 ,n2063);
    or g704(n2229 ,n1910 ,n2083);
    or g705(n2228 ,n1802 ,n2108);
    or g706(n2227 ,n2094 ,n1956);
    or g707(n2226 ,n1797 ,n2142);
    or g708(n2225 ,n1798 ,n2060);
    or g709(n2224 ,n1917 ,n2059);
    or g710(n2223 ,n2163 ,n1934);
    or g711(n2222 ,n1700 ,n2165);
    or g712(n2221 ,n1701 ,n2164);
    or g713(n2220 ,n1699 ,n2166);
    or g714(n2219 ,n1852 ,n2057);
    or g715(n2218 ,n1851 ,n2055);
    or g716(n2217 ,n1853 ,n2056);
    or g717(n2216 ,n1850 ,n2054);
    or g718(n2215 ,n1849 ,n2053);
    or g719(n2214 ,n1848 ,n2052);
    or g720(n2213 ,n1924 ,n2050);
    or g721(n2212 ,n1846 ,n2048);
    or g722(n2211 ,n1845 ,n2047);
    or g723(n2210 ,n1843 ,n2046);
    or g724(n2209 ,n1842 ,n2045);
    or g725(n2208 ,n1840 ,n2044);
    or g726(n2207 ,n1923 ,n2042);
    or g727(n2206 ,n1841 ,n2043);
    or g728(n2205 ,n1838 ,n2040);
    or g729(n2204 ,n1837 ,n2039);
    or g730(n2203 ,n1836 ,n2038);
    or g731(n2202 ,n1835 ,n2037);
    or g732(n2201 ,n1834 ,n2036);
    or g733(n2200 ,n1833 ,n2035);
    or g734(n2199 ,n1922 ,n2034);
    or g735(n2198 ,n1831 ,n2031);
    or g736(n2197 ,n1830 ,n2030);
    or g737(n2196 ,n1829 ,n2029);
    or g738(n2195 ,n1828 ,n2028);
    or g739(n2194 ,n1826 ,n2026);
    or g740(n2193 ,n1827 ,n2027);
    or g741(n2192 ,n1921 ,n2025);
    or g742(n2191 ,n1824 ,n2023);
    or g743(n2190 ,n1823 ,n2021);
    or g744(n2189 ,n1822 ,n2022);
    or g745(n2188 ,n1821 ,n2020);
    or g746(n2187 ,n1928 ,n2102);
    or g747(n2186 ,n1820 ,n2019);
    or g748(n2185 ,n1819 ,n2018);
    or g749(n2184 ,n1920 ,n2017);
    or g750(n2183 ,n1816 ,n2014);
    or g751(n2182 ,n1814 ,n2012);
    or g752(n2181 ,n1813 ,n2011);
    or g753(n2180 ,n1815 ,n2013);
    or g754(n2179 ,n1812 ,n2010);
    or g755(n2178 ,n1811 ,n2009);
    or g756(n2177 ,n1919 ,n2008);
    or g757(n2176 ,n1809 ,n2006);
    or g758(n2175 ,n1808 ,n2005);
    or g759(n2174 ,n1807 ,n2004);
    or g760(n2173 ,n1806 ,n2003);
    or g761(n2172 ,n1805 ,n2002);
    or g762(n2171 ,n1803 ,n2001);
    or g763(n2170 ,n1918 ,n2000);
    nor g764(n2169 ,n553 ,n1968);
    nor g765(n2168 ,n598 ,n1873);
    nor g766(n2167 ,n580 ,n1969);
    nor g767(n2166 ,n362 ,n1876);
    nor g768(n2165 ,n385 ,n1876);
    nor g769(n2164 ,n392 ,n1876);
    nor g770(n2163 ,n433 ,n1874);
    nor g771(n2162 ,n231 ,n1874);
    nor g772(n2161 ,n226 ,n1874);
    nor g773(n2160 ,n227 ,n1874);
    nor g774(n2159 ,n581 ,n1869);
    nor g775(n2158 ,n269 ,n1869);
    nor g776(n2157 ,n495 ,n1869);
    nor g777(n2156 ,n524 ,n1869);
    nor g778(n2155 ,n545 ,n1869);
    nor g779(n2154 ,n494 ,n1869);
    nor g780(n2153 ,n440 ,n1967);
    nor g781(n2152 ,n307 ,n1869);
    nor g782(n2151 ,n479 ,n1860);
    nor g783(n2150 ,n324 ,n1860);
    nor g784(n2149 ,n478 ,n1860);
    nor g785(n2148 ,n512 ,n1860);
    nor g786(n2147 ,n563 ,n1860);
    nor g787(n2146 ,n474 ,n1860);
    nor g788(n2145 ,n312 ,n1860);
    nor g789(n2144 ,n313 ,n1860);
    nor g790(n2143 ,n472 ,n1861);
    nor g791(n2142 ,n544 ,n1873);
    nor g792(n2141 ,n263 ,n1861);
    nor g793(n2140 ,n302 ,n1861);
    nor g794(n2139 ,n590 ,n1969);
    nor g795(n2138 ,n338 ,n1861);
    nor g796(n2137 ,n259 ,n1861);
    nor g797(n2136 ,n273 ,n1861);
    nor g798(n2135 ,n448 ,n1861);
    nor g799(n2134 ,n275 ,n1861);
    nor g800(n2133 ,n520 ,n1865);
    nor g801(n2132 ,n586 ,n1865);
    nor g802(n2131 ,n349 ,n1865);
    nor g803(n2130 ,n530 ,n1865);
    nor g804(n2129 ,n294 ,n1865);
    nor g805(n2128 ,n276 ,n1865);
    nor g806(n2127 ,n589 ,n1865);
    nor g807(n2126 ,n317 ,n1865);
    nor g808(n2125 ,n497 ,n1862);
    nor g809(n2124 ,n291 ,n1862);
    nor g810(n2123 ,n525 ,n1968);
    nor g811(n2122 ,n503 ,n1862);
    nor g812(n2121 ,n306 ,n1969);
    nor g813(n2120 ,n235 ,n1862);
    nor g814(n2119 ,n242 ,n1862);
    nor g815(n2118 ,n516 ,n1862);
    nor g816(n2117 ,n508 ,n1862);
    nor g817(n2116 ,n454 ,n1967);
    nor g818(n2115 ,n517 ,n1864);
    nor g819(n2114 ,n579 ,n1967);
    nor g820(n2113 ,n555 ,n1863);
    nor g821(n2112 ,n353 ,n1968);
    nor g822(n2111 ,n542 ,n1863);
    nor g823(n2110 ,n350 ,n1863);
    nor g824(n2109 ,n339 ,n1967);
    nor g825(n2108 ,n237 ,n1873);
    nor g826(n2107 ,n552 ,n1863);
    nor g827(n2106 ,n283 ,n1863);
    nor g828(n2105 ,n461 ,n1968);
    nor g829(n2104 ,n582 ,n1969);
    nor g830(n2103 ,n304 ,n1863);
    nor g831(n2102 ,n526 ,n1863);
    nor g832(n2101 ,n285 ,n1859);
    nor g833(n2100 ,n333 ,n1859);
    nor g834(n2099 ,n240 ,n1968);
    nor g835(n2098 ,n327 ,n1859);
    nor g836(n2097 ,n345 ,n1864);
    nor g837(n2096 ,n331 ,n1969);
    nor g838(n2095 ,n329 ,n1859);
    nor g839(n2094 ,n278 ,n1969);
    nor g840(n2093 ,n551 ,n1859);
    nor g841(n2092 ,n352 ,n1968);
    nor g842(n2091 ,n515 ,n1859);
    nor g843(n2090 ,n578 ,n1969);
    nor g844(n2089 ,n564 ,n1859);
    nor g845(n2088 ,n321 ,n1967);
    nor g846(n2087 ,n504 ,n1967);
    nor g847(n2086 ,n575 ,n1864);
    nor g848(n2085 ,n556 ,n1864);
    nor g849(n2084 ,n298 ,n1968);
    nor g850(n2083 ,n450 ,n1864);
    nor g851(n2082 ,n279 ,n1864);
    nor g852(n2081 ,n340 ,n1859);
    nor g853(n2080 ,n477 ,n1864);
    nor g854(n2079 ,n289 ,n1862);
    nor g855(n2078 ,n522 ,n1864);
    nor g856(n2077 ,n539 ,n1968);
    or g857(n2064 ,n1961 ,n1793);
    nor g858(n2063 ,n559 ,n1873);
    nor g859(n2062 ,n443 ,n1873);
    nor g860(n2061 ,n260 ,n1967);
    nor g861(n2060 ,n320 ,n1873);
    nor g862(n2059 ,n583 ,n1873);
    nor g863(n2058 ,n567 ,n1866);
    nor g864(n2057 ,n561 ,n1866);
    nor g865(n2056 ,n587 ,n1866);
    nor g866(n2055 ,n261 ,n1866);
    nor g867(n2054 ,n249 ,n1866);
    nor g868(n2053 ,n510 ,n1866);
    nor g869(n2052 ,n305 ,n1866);
    nor g870(n2051 ,n493 ,n1969);
    nor g871(n2050 ,n234 ,n1866);
    nor g872(n2049 ,n347 ,n1868);
    nor g873(n2048 ,n233 ,n1868);
    nor g874(n2047 ,n300 ,n1868);
    nor g875(n2046 ,n456 ,n1868);
    nor g876(n2045 ,n244 ,n1868);
    nor g877(n2044 ,n505 ,n1868);
    nor g878(n2043 ,n513 ,n1868);
    nor g879(n2042 ,n466 ,n1868);
    nor g880(n2041 ,n546 ,n1867);
    nor g881(n2040 ,n270 ,n1867);
    nor g882(n2039 ,n292 ,n1867);
    nor g883(n2038 ,n355 ,n1867);
    nor g884(n2037 ,n585 ,n1867);
    nor g885(n2036 ,n458 ,n1867);
    nor g886(n2035 ,n336 ,n1867);
    nor g887(n2034 ,n481 ,n1867);
    nor g888(n2033 ,n441 ,n1967);
    nor g889(n2032 ,n566 ,n1858);
    nor g890(n2031 ,n490 ,n1858);
    nor g891(n2030 ,n550 ,n1858);
    nor g892(n2029 ,n451 ,n1858);
    nor g893(n2028 ,n287 ,n1858);
    nor g894(n2027 ,n284 ,n1858);
    nor g895(n2026 ,n264 ,n1858);
    nor g896(n2025 ,n509 ,n1858);
    nor g897(n2024 ,n488 ,n1872);
    nor g898(n2023 ,n319 ,n1872);
    nor g899(n2022 ,n314 ,n1872);
    nor g900(n2021 ,n281 ,n1872);
    nor g901(n2020 ,n571 ,n1872);
    nor g902(n2019 ,n492 ,n1872);
    nor g903(n2018 ,n251 ,n1872);
    nor g904(n2017 ,n444 ,n1872);
    nor g905(n2016 ,n527 ,n1863);
    nor g906(n2015 ,n475 ,n1871);
    nor g907(n2014 ,n262 ,n1871);
    nor g908(n2013 ,n265 ,n1871);
    nor g909(n2012 ,n344 ,n1871);
    nor g910(n2011 ,n521 ,n1871);
    nor g911(n2010 ,n301 ,n1871);
    nor g912(n2009 ,n247 ,n1871);
    nor g913(n2008 ,n588 ,n1871);
    nor g914(n2007 ,n463 ,n1870);
    nor g915(n2006 ,n507 ,n1870);
    nor g916(n2005 ,n351 ,n1870);
    nor g917(n2004 ,n518 ,n1870);
    nor g918(n2003 ,n572 ,n1870);
    nor g919(n2002 ,n560 ,n1870);
    nor g920(n2001 ,n342 ,n1870);
    nor g921(n2000 ,n238 ,n1870);
    nor g922(n1999 ,n256 ,n1869);
    nor g923(n1998 ,n412 ,n1874);
    nor g924(n1997 ,n584 ,n1873);
    or g925(n1996 ,n195 ,n1810);
    or g926(n1995 ,n201 ,n1817);
    or g927(n1994 ,n199 ,n1825);
    or g928(n1993 ,n202 ,n1832);
    or g929(n1992 ,n194 ,n1839);
    or g930(n1991 ,n199 ,n1847);
    or g931(n1990 ,n194 ,n1854);
    or g932(n1989 ,n195 ,n1796);
    or g933(n1988 ,n199 ,n1965);
    or g934(n1987 ,n201 ,n1937);
    or g935(n1986 ,n194 ,n1877);
    or g936(n1985 ,n1740 ,n1933);
    or g937(n1984 ,n1960 ,n1777);
    or g938(n1983 ,n1959 ,n1857);
    or g939(n1982 ,n1958 ,n1778);
    or g940(n1981 ,n1940 ,n1782);
    or g941(n1980 ,n1472 ,n1785);
    or g942(n1979 ,n201 ,n1916);
    or g943(n1978 ,n194 ,n1908);
    or g944(n1977 ,n195 ,n1901);
    or g945(n1976 ,n195 ,n1894);
    nor g946(n1975 ,n198 ,n1779);
    nor g947(n1974 ,n196 ,n1780);
    nor g948(n1973 ,n196 ,n1781);
    or g949(n1972 ,n201 ,n1888);
    or g950(n2076 ,n643 ,n1970);
    or g951(n2075 ,n614 ,n1970);
    or g952(n2074 ,n614 ,n1875);
    or g953(n2073 ,n648 ,n1875);
    or g954(n2072 ,n648 ,n1971);
    or g955(n2071 ,n646 ,n1875);
    or g956(n2070 ,n614 ,n1971);
    or g957(n2069 ,n643 ,n1875);
    or g958(n2068 ,n643 ,n1971);
    or g959(n2067 ,n646 ,n1970);
    or g960(n2066 ,n648 ,n1970);
    or g961(n2065 ,n646 ,n1971);
    nor g962(n1966 ,n404 ,n1766);
    nor g963(n1965 ,n205 ,n1772);
    nor g964(n1964 ,n404 ,n1772);
    nor g965(n1963 ,n403 ,n1774);
    nor g966(n1962 ,n206 ,n1772);
    nor g967(n1961 ,n428 ,n1735);
    nor g968(n1960 ,n436 ,n1735);
    nor g969(n1959 ,n427 ,n1735);
    nor g970(n1958 ,n437 ,n1735);
    nor g971(n1957 ,n335 ,n1733);
    nor g972(n1956 ,n257 ,n1733);
    nor g973(n1955 ,n328 ,n1732);
    nor g974(n1954 ,n246 ,n1733);
    nor g975(n1953 ,n499 ,n1732);
    nor g976(n1952 ,n299 ,n1733);
    nor g977(n1951 ,n330 ,n1732);
    nor g978(n1950 ,n267 ,n1733);
    nor g979(n1949 ,n252 ,n1732);
    nor g980(n1948 ,n489 ,n1733);
    nor g981(n1947 ,n574 ,n1733);
    nor g982(n1946 ,n293 ,n1732);
    nor g983(n1945 ,n348 ,n1732);
    nor g984(n1944 ,n462 ,n1733);
    nor g985(n1943 ,n533 ,n1732);
    nor g986(n1942 ,n245 ,n1732);
    nor g987(n1941 ,n405 ,n1768);
    nor g988(n1940 ,n222 ,n1735);
    nor g989(n1939 ,n204 ,n1768);
    or g990(n1938 ,n1158 ,n1719);
    nor g991(n1937 ,n205 ,n1768);
    nor g992(n1936 ,n405 ,n1766);
    nor g993(n1935 ,n206 ,n1768);
    nor g994(n1934 ,n626 ,n1739);
    or g995(n1933 ,n1720 ,n1681);
    nor g996(n1932 ,n406 ,n1764);
    nor g997(n1931 ,n406 ,n1762);
    nor g998(n1930 ,n406 ,n1776);
    nor g999(n1929 ,n406 ,n1774);
    nor g1000(n1928 ,n406 ,n1768);
    nor g1001(n1927 ,n406 ,n1766);
    nor g1002(n1926 ,n406 ,n1772);
    nor g1003(n1925 ,n406 ,n1770);
    nor g1004(n1924 ,n406 ,n1760);
    nor g1005(n1923 ,n406 ,n1758);
    nor g1006(n1922 ,n406 ,n1756);
    nor g1007(n1921 ,n406 ,n1754);
    nor g1008(n1920 ,n406 ,n1727);
    nor g1009(n1919 ,n406 ,n1731);
    nor g1010(n1918 ,n406 ,n1729);
    nor g1011(n1917 ,n406 ,n1751);
    nor g1012(n1916 ,n205 ,n1764);
    nor g1013(n1915 ,n204 ,n1764);
    nor g1014(n1914 ,n206 ,n1764);
    nor g1015(n1913 ,n405 ,n1764);
    nor g1016(n1912 ,n404 ,n1764);
    nor g1017(n1911 ,n402 ,n1764);
    nor g1018(n1910 ,n405 ,n1772);
    nor g1019(n1909 ,n403 ,n1764);
    nor g1020(n1908 ,n205 ,n1762);
    nor g1021(n1907 ,n204 ,n1762);
    nor g1022(n1906 ,n206 ,n1762);
    nor g1023(n1905 ,n405 ,n1762);
    nor g1024(n1904 ,n404 ,n1762);
    nor g1025(n1903 ,n402 ,n1762);
    nor g1026(n1902 ,n403 ,n1762);
    nor g1027(n1901 ,n205 ,n1776);
    nor g1028(n1900 ,n204 ,n1776);
    nor g1029(n1899 ,n206 ,n1776);
    nor g1030(n1898 ,n405 ,n1776);
    nor g1031(n1897 ,n404 ,n1776);
    nor g1032(n1896 ,n402 ,n1776);
    nor g1033(n1895 ,n403 ,n1776);
    nor g1034(n1894 ,n205 ,n1774);
    nor g1035(n1893 ,n204 ,n1774);
    nor g1036(n1892 ,n204 ,n1772);
    nor g1037(n1891 ,n404 ,n1774);
    nor g1038(n1890 ,n402 ,n1766);
    nor g1039(n1889 ,n206 ,n1774);
    nor g1040(n1888 ,n205 ,n1770);
    nor g1041(n1887 ,n204 ,n1770);
    nor g1042(n1886 ,n405 ,n1770);
    nor g1043(n1885 ,n404 ,n1770);
    nor g1044(n1884 ,n403 ,n1772);
    nor g1045(n1883 ,n402 ,n1770);
    nor g1046(n1882 ,n403 ,n1770);
    nor g1047(n1881 ,n206 ,n1770);
    nor g1048(n1880 ,n402 ,n1774);
    nor g1049(n1879 ,n402 ,n1772);
    nor g1050(n1878 ,n402 ,n1768);
    nor g1051(n1877 ,n205 ,n1766);
    or g1052(n1971 ,n217 ,n1737);
    or g1053(n1970 ,n418 ,n1712);
    or g1054(n1969 ,n648 ,n1736);
    or g1055(n1968 ,n646 ,n1736);
    or g1056(n1967 ,n614 ,n1736);
    or g1057(n1857 ,n772 ,n1746);
    nor g1058(n1856 ,n403 ,n1766);
    nor g1059(n1855 ,n206 ,n1766);
    nor g1060(n1854 ,n205 ,n1760);
    nor g1061(n1853 ,n204 ,n1760);
    nor g1062(n1852 ,n206 ,n1760);
    nor g1063(n1851 ,n405 ,n1760);
    nor g1064(n1850 ,n404 ,n1760);
    nor g1065(n1849 ,n402 ,n1760);
    nor g1066(n1848 ,n403 ,n1760);
    nor g1067(n1847 ,n205 ,n1758);
    nor g1068(n1846 ,n204 ,n1758);
    nor g1069(n1845 ,n206 ,n1758);
    nor g1070(n1844 ,n204 ,n1766);
    nor g1071(n1843 ,n405 ,n1758);
    nor g1072(n1842 ,n404 ,n1758);
    nor g1073(n1841 ,n403 ,n1758);
    nor g1074(n1840 ,n402 ,n1758);
    nor g1075(n1839 ,n205 ,n1756);
    nor g1076(n1838 ,n204 ,n1756);
    nor g1077(n1837 ,n206 ,n1756);
    nor g1078(n1836 ,n405 ,n1756);
    nor g1079(n1835 ,n404 ,n1756);
    nor g1080(n1834 ,n402 ,n1756);
    nor g1081(n1833 ,n403 ,n1756);
    nor g1082(n1832 ,n205 ,n1754);
    nor g1083(n1831 ,n204 ,n1754);
    nor g1084(n1830 ,n206 ,n1754);
    nor g1085(n1829 ,n405 ,n1754);
    nor g1086(n1828 ,n404 ,n1754);
    nor g1087(n1827 ,n402 ,n1754);
    nor g1088(n1826 ,n403 ,n1754);
    nor g1089(n1825 ,n205 ,n1727);
    nor g1090(n1824 ,n204 ,n1727);
    nor g1091(n1823 ,n206 ,n1727);
    nor g1092(n1822 ,n405 ,n1727);
    nor g1093(n1821 ,n404 ,n1727);
    nor g1094(n1820 ,n402 ,n1727);
    nor g1095(n1819 ,n403 ,n1727);
    nor g1096(n1818 ,n403 ,n1768);
    nor g1097(n1817 ,n205 ,n1731);
    nor g1098(n1816 ,n204 ,n1731);
    nor g1099(n1815 ,n206 ,n1731);
    nor g1100(n1814 ,n405 ,n1731);
    nor g1101(n1813 ,n404 ,n1731);
    nor g1102(n1812 ,n402 ,n1731);
    nor g1103(n1811 ,n403 ,n1731);
    nor g1104(n1810 ,n205 ,n1729);
    nor g1105(n1809 ,n204 ,n1729);
    nor g1106(n1808 ,n206 ,n1729);
    nor g1107(n1807 ,n405 ,n1729);
    nor g1108(n1806 ,n404 ,n1729);
    nor g1109(n1805 ,n402 ,n1729);
    nor g1110(n1804 ,n404 ,n1768);
    nor g1111(n1803 ,n403 ,n1729);
    nor g1112(n1802 ,n405 ,n1751);
    nor g1113(n1801 ,n204 ,n1751);
    nor g1114(n1800 ,n206 ,n1751);
    nor g1115(n1799 ,n402 ,n1751);
    nor g1116(n1798 ,n403 ,n1751);
    nor g1117(n1797 ,n404 ,n1751);
    nor g1118(n1796 ,n205 ,n1751);
    or g1119(n1795 ,n1088 ,n1718);
    or g1120(n1794 ,n1080 ,n1714);
    nor g1121(n1793 ,n627 ,n1734);
    or g1122(n1792 ,n1008 ,n1715);
    nor g1123(n1791 ,n405 ,n1774);
    or g1124(n1790 ,n1055 ,n1725);
    or g1125(n1789 ,n1040 ,n1711);
    or g1126(n1788 ,n1010 ,n1710);
    or g1127(n1787 ,n1075 ,n1709);
    or g1128(n1786 ,n1644 ,n1742);
    or g1129(n1785 ,n1590 ,n1722);
    or g1130(n1784 ,n1743 ,n1741);
    nor g1131(n1783 ,n197 ,n1724);
    or g1132(n1782 ,n771 ,n1750);
    nor g1133(n1781 ,n1703 ,n1748);
    nor g1134(n1780 ,n1704 ,n1749);
    nor g1135(n1779 ,n1702 ,n1744);
    or g1136(n1778 ,n770 ,n1745);
    or g1137(n1777 ,n769 ,n1747);
    or g1138(n1876 ,n1624 ,n1752);
    or g1139(n1875 ,n58[0] ,n1737);
    or g1140(n1874 ,n195 ,n1738);
    or g1141(n1873 ,n199 ,n1752);
    or g1142(n1872 ,n202 ,n1726);
    or g1143(n1871 ,n200 ,n1730);
    or g1144(n1870 ,n201 ,n1728);
    or g1145(n1869 ,n202 ,n1763);
    or g1146(n1868 ,n200 ,n1757);
    or g1147(n1867 ,n195 ,n1755);
    or g1148(n1866 ,n200 ,n1759);
    or g1149(n1865 ,n199 ,n1773);
    or g1150(n1864 ,n202 ,n1771);
    or g1151(n1863 ,n200 ,n1767);
    or g1152(n1862 ,n200 ,n1769);
    or g1153(n1861 ,n200 ,n1775);
    or g1154(n1860 ,n202 ,n1761);
    or g1155(n1859 ,n201 ,n1765);
    or g1156(n1858 ,n199 ,n1753);
    not g1157(n1776 ,n1775);
    not g1158(n1774 ,n1773);
    not g1159(n1772 ,n1771);
    not g1160(n1770 ,n1769);
    not g1161(n1768 ,n1767);
    not g1162(n1766 ,n1765);
    not g1163(n1764 ,n1763);
    not g1164(n1762 ,n1761);
    not g1165(n1760 ,n1759);
    not g1166(n1758 ,n1757);
    not g1167(n1756 ,n1755);
    not g1168(n1754 ,n1753);
    not g1169(n1751 ,n1752);
    nor g1170(n1750 ,n361 ,n1689);
    nor g1171(n1749 ,n367 ,n185);
    nor g1172(n1748 ,n370 ,n185);
    nor g1173(n1747 ,n376 ,n1689);
    nor g1174(n1746 ,n384 ,n1689);
    nor g1175(n1745 ,n382 ,n1689);
    nor g1176(n1744 ,n393 ,n185);
    nor g1177(n1743 ,n407 ,n1692);
    nor g1178(n1742 ,n203 ,n1692);
    nor g1179(n1741 ,n1139 ,n1674);
    or g1180(n1740 ,n1635 ,n1679);
    nor g1181(n1775 ,n615 ,n1707);
    nor g1182(n1773 ,n649 ,n1708);
    nor g1183(n1771 ,n644 ,n1708);
    nor g1184(n1769 ,n649 ,n1707);
    nor g1185(n1767 ,n650 ,n1708);
    nor g1186(n1765 ,n650 ,n1707);
    nor g1187(n1763 ,n644 ,n1691);
    nor g1188(n1761 ,n615 ,n1708);
    nor g1189(n1759 ,n615 ,n1690);
    nor g1190(n1757 ,n615 ,n1691);
    nor g1191(n1755 ,n649 ,n1690);
    nor g1192(n1753 ,n649 ,n1691);
    nor g1193(n1752 ,n644 ,n1707);
    not g1194(n1739 ,n1738);
    not g1195(n1735 ,n1734);
    not g1196(n1731 ,n1730);
    not g1197(n1729 ,n1728);
    not g1198(n1727 ,n1726);
    or g1199(n1725 ,n996 ,n1686);
    xnor g1200(n1724 ,n1670 ,n58[0]);
    or g1201(n1723 ,n1664 ,n1697);
    nor g1202(n1722 ,n401 ,n1692);
    or g1203(n1721 ,n1656 ,n1694);
    or g1204(n1720 ,n1696 ,n1695);
    or g1205(n1719 ,n202 ,n1687);
    or g1206(n1718 ,n1002 ,n1676);
    or g1207(n1717 ,n1646 ,n1698);
    or g1208(n1716 ,n1658 ,n1680);
    or g1209(n1715 ,n1001 ,n1688);
    or g1210(n1714 ,n1000 ,n1684);
    or g1211(n1713 ,n1659 ,n1706);
    or g1212(n1712 ,n58[0] ,n1689);
    or g1213(n1711 ,n995 ,n1683);
    or g1214(n1710 ,n999 ,n1682);
    or g1215(n1709 ,n997 ,n1705);
    nor g1216(n1738 ,n605 ,n1672);
    or g1217(n1737 ,n58[1] ,n1689);
    or g1218(n1736 ,n656 ,n1689);
    nor g1219(n1734 ,n737 ,n1693);
    or g1220(n1733 ,n1521 ,n1693);
    or g1221(n1732 ,n680 ,n1689);
    nor g1222(n1730 ,n650 ,n1691);
    nor g1223(n1728 ,n644 ,n1690);
    nor g1224(n1726 ,n650 ,n1690);
    nor g1225(n1706 ,n379 ,n187);
    or g1226(n1705 ,n1490 ,n1655);
    nor g1227(n1704 ,n415 ,n1670);
    nor g1228(n1703 ,n218 ,n1670);
    nor g1229(n1702 ,n418 ,n1670);
    nor g1230(n1701 ,n410 ,n1645);
    nor g1231(n1700 ,n411 ,n1645);
    nor g1232(n1699 ,n414 ,n1645);
    nor g1233(n1698 ,n221 ,n1645);
    nor g1234(n1697 ,n381 ,n187);
    nor g1235(n1696 ,n364 ,n1657);
    nor g1236(n1695 ,n386 ,n1637);
    nor g1237(n1694 ,n390 ,n187);
    or g1238(n1708 ,n410 ,n1647);
    or g1239(n1707 ,n410 ,n186);
    or g1240(n1688 ,n1465 ,n1652);
    or g1241(n1687 ,n1480 ,n1668);
    or g1242(n1686 ,n1477 ,n1654);
    nor g1243(n1685 ,n1529 ,n1626);
    or g1244(n1684 ,n1482 ,n1651);
    or g1245(n1683 ,n1470 ,n1643);
    or g1246(n1682 ,n1467 ,n1642);
    or g1247(n1681 ,n1666 ,n1665);
    nor g1248(n1680 ,n672 ,n1638);
    or g1249(n1679 ,n1667 ,n1650);
    or g1250(n1678 ,n747 ,n1660);
    or g1251(n1677 ,n748 ,n1661);
    or g1252(n1676 ,n1487 ,n1653);
    nor g1253(n1675 ,n196 ,n1636);
    or g1254(n1674 ,n199 ,n1648);
    or g1255(n1673 ,n749 ,n1662);
    or g1256(n1672 ,n18[1] ,n1634);
    or g1257(n1671 ,n753 ,n1663);
    or g1258(n1693 ,n201 ,n1670);
    or g1259(n1692 ,n195 ,n1649);
    or g1260(n1691 ,n40[3] ,n186);
    or g1261(n1690 ,n40[3] ,n1647);
    or g1262(n1689 ,n202 ,n1669);
    not g1263(n1669 ,n1670);
    or g1264(n1668 ,n1147 ,n1583);
    nor g1265(n1667 ,n375 ,n1617);
    nor g1266(n1666 ,n395 ,n1619);
    nor g1267(n1665 ,n377 ,n1620);
    nor g1268(n1664 ,n438 ,n1606);
    nor g1269(n1663 ,n274 ,n1624);
    nor g1270(n1662 ,n250 ,n1624);
    nor g1271(n1661 ,n243 ,n1624);
    nor g1272(n1660 ,n241 ,n1624);
    nor g1273(n1659 ,n220 ,n1606);
    nor g1274(n1658 ,n409 ,n1606);
    or g1275(n1657 ,n216 ,n1625);
    nor g1276(n1656 ,n216 ,n1606);
    or g1277(n1655 ,n1186 ,n1589);
    or g1278(n1654 ,n1131 ,n1584);
    or g1279(n1653 ,n1165 ,n1588);
    or g1280(n1652 ,n1152 ,n1587);
    or g1281(n1651 ,n1161 ,n1586);
    nor g1282(n1650 ,n365 ,n1618);
    nor g1283(n1670 ,n633 ,n1577);
    not g1284(n1649 ,n1648);
    not g1285(n1647 ,n1646);
    nor g1286(n1644 ,n196 ,n1591);
    or g1287(n1643 ,n1132 ,n1582);
    or g1288(n1642 ,n1176 ,n1581);
    or g1289(n1641 ,n654 ,n1574);
    or g1290(n1640 ,n1540 ,n1578);
    or g1291(n1639 ,n1528 ,n1585);
    or g1292(n1638 ,n21[0] ,n1605);
    or g1293(n1637 ,n21[2] ,n1625);
    nor g1294(n1636 ,n11[3] ,n1615);
    or g1295(n1635 ,n1607 ,n1613);
    nor g1296(n1634 ,n618 ,n1616);
    or g1297(n1633 ,n1604 ,n1603);
    or g1298(n1632 ,n1601 ,n1602);
    or g1299(n1631 ,n1600 ,n1599);
    or g1300(n1630 ,n1597 ,n1598);
    or g1301(n1629 ,n1596 ,n1595);
    or g1302(n1628 ,n1593 ,n1594);
    or g1303(n1627 ,n1621 ,n1592);
    or g1304(n1626 ,n1518 ,n1573);
    nor g1305(n1648 ,n1579 ,n1580);
    nor g1306(n1646 ,n40[0] ,n1624);
    or g1307(n1645 ,n198 ,n1623);
    not g1308(n1624 ,n1623);
    nor g1309(n1622 ,n489 ,n1563);
    nor g1310(n1621 ,n406 ,n1564);
    or g1311(n1620 ,n621 ,n1566);
    or g1312(n1619 ,n621 ,n1572);
    or g1313(n1618 ,n653 ,n1566);
    or g1314(n1617 ,n653 ,n1572);
    nor g1315(n1616 ,n203 ,n1569);
    nor g1316(n1615 ,n412 ,n1531);
    nor g1317(n1614 ,n299 ,n1563);
    nor g1318(n1613 ,n257 ,n1563);
    nor g1319(n1612 ,n574 ,n1563);
    nor g1320(n1611 ,n246 ,n1563);
    nor g1321(n1610 ,n335 ,n1563);
    nor g1322(n1609 ,n267 ,n1563);
    nor g1323(n1608 ,n462 ,n1563);
    nor g1324(n1607 ,n387 ,n1536);
    or g1325(n1625 ,n409 ,n1566);
    nor g1326(n1623 ,n673 ,n1569);
    nor g1327(n1604 ,n204 ,n1564);
    nor g1328(n1603 ,n205 ,n1565);
    nor g1329(n1602 ,n204 ,n1565);
    nor g1330(n1601 ,n206 ,n1564);
    nor g1331(n1600 ,n405 ,n1564);
    nor g1332(n1599 ,n206 ,n1565);
    nor g1333(n1598 ,n405 ,n1565);
    nor g1334(n1597 ,n404 ,n1564);
    nor g1335(n1596 ,n402 ,n1564);
    nor g1336(n1595 ,n404 ,n1565);
    nor g1337(n1594 ,n402 ,n1565);
    nor g1338(n1593 ,n403 ,n1564);
    nor g1339(n1592 ,n403 ,n1565);
    nor g1340(n1591 ,n1463 ,n1542);
    nor g1341(n1590 ,n197 ,n1556);
    or g1342(n1589 ,n1067 ,n1530);
    or g1343(n1588 ,n1109 ,n1532);
    or g1344(n1587 ,n1092 ,n1533);
    or g1345(n1586 ,n1069 ,n1534);
    or g1346(n1585 ,n1231 ,n1541);
    or g1347(n1584 ,n1046 ,n1535);
    or g1348(n1583 ,n1043 ,n1537);
    or g1349(n1582 ,n1019 ,n1538);
    or g1350(n1581 ,n1110 ,n1539);
    nor g1351(n1580 ,n401 ,n1555);
    nor g1352(n1579 ,n18[1] ,n1554);
    or g1353(n1578 ,n198 ,n1527);
    or g1354(n1577 ,n18[1] ,n1557);
    or g1355(n1576 ,n655 ,n1571);
    or g1356(n1575 ,n657 ,n1570);
    or g1357(n1574 ,n1571 ,n1570);
    nor g1358(n1573 ,n18[1] ,n1553);
    or g1359(n1606 ,n195 ,n1567);
    or g1360(n1605 ,n201 ,n1568);
    not g1361(n1568 ,n1567);
    or g1362(n1562 ,n708 ,n1493);
    or g1363(n1561 ,n724 ,n1494);
    or g1364(n1560 ,n720 ,n1495);
    or g1365(n1559 ,n722 ,n1497);
    or g1366(n1558 ,n704 ,n1496);
    nor g1367(n1557 ,n1226 ,n1459);
    or g1368(n1556 ,n660 ,n1421);
    nor g1369(n1555 ,n1461 ,n1422);
    nor g1370(n1554 ,n662 ,n1525);
    nor g1371(n1553 ,n1226 ,n1522);
    or g1372(n1552 ,n717 ,n1492);
    or g1373(n1551 ,n721 ,n1501);
    or g1374(n1550 ,n710 ,n1503);
    or g1375(n1549 ,n718 ,n1500);
    or g1376(n1548 ,n715 ,n1499);
    or g1377(n1547 ,n723 ,n1504);
    or g1378(n1546 ,n725 ,n1498);
    or g1379(n1545 ,n709 ,n1505);
    or g1380(n1544 ,n714 ,n1506);
    or g1381(n1543 ,n719 ,n1507);
    nor g1382(n1542 ,n18[1] ,n1526);
    nor g1383(n1541 ,n14 ,n1437);
    nor g1384(n1540 ,n205 ,n1516);
    or g1385(n1539 ,n1466 ,n1464);
    or g1386(n1538 ,n1515 ,n1468);
    or g1387(n1537 ,n1473 ,n1471);
    or g1388(n1536 ,n658 ,n1519);
    or g1389(n1535 ,n1475 ,n1474);
    or g1390(n1534 ,n1481 ,n1479);
    or g1391(n1533 ,n1484 ,n1483);
    or g1392(n1532 ,n1486 ,n1485);
    or g1393(n1531 ,n617 ,n1523);
    or g1394(n1530 ,n1489 ,n1488);
    or g1395(n1529 ,n562 ,n1521);
    nor g1396(n1528 ,n421 ,n1436);
    nor g1397(n1527 ,n229 ,n1517);
    or g1398(n1572 ,n220 ,n1519);
    nor g1399(n1571 ,n629 ,n1524);
    nor g1400(n1570 ,n669 ,n1524);
    or g1401(n1569 ,n20[4] ,n1523);
    nor g1402(n1567 ,n620 ,n1424);
    or g1403(n1566 ,n21[1] ,n1519);
    or g1404(n1565 ,n194 ,n1517);
    or g1405(n1564 ,n199 ,n1516);
    or g1406(n1563 ,n201 ,n1520);
    not g1407(n1526 ,n1525);
    not g1408(n1523 ,n1522);
    not g1409(n1520 ,n1521);
    not g1410(n1519 ,n1518);
    not g1411(n1517 ,n1516);
    or g1412(n1515 ,n1130 ,n1127);
    or g1413(n1514 ,n915 ,n1312);
    or g1414(n1513 ,n907 ,n1313);
    or g1415(n1512 ,n888 ,n1315);
    or g1416(n1511 ,n868 ,n1317);
    or g1417(n1510 ,n863 ,n1318);
    or g1418(n1509 ,n945 ,n1320);
    or g1419(n1508 ,n859 ,n1321);
    nor g1420(n1507 ,n374 ,n192);
    nor g1421(n1506 ,n389 ,n190);
    nor g1422(n1505 ,n368 ,n189);
    nor g1423(n1504 ,n398 ,n188);
    nor g1424(n1503 ,n363 ,n193);
    or g1425(n1502 ,n931 ,n1322);
    nor g1426(n1501 ,n397 ,n190);
    nor g1427(n1500 ,n372 ,n188);
    nor g1428(n1499 ,n399 ,n189);
    nor g1429(n1498 ,n383 ,n191);
    nor g1430(n1497 ,n378 ,n193);
    nor g1431(n1496 ,n369 ,n192);
    nor g1432(n1495 ,n373 ,n191);
    nor g1433(n1494 ,n394 ,n192);
    nor g1434(n1493 ,n366 ,n191);
    nor g1435(n1492 ,n391 ,n191);
    or g1436(n1491 ,n911 ,n1324);
    or g1437(n1490 ,n1170 ,n1190);
    or g1438(n1489 ,n1181 ,n1163);
    or g1439(n1488 ,n1187 ,n1154);
    or g1440(n1487 ,n1185 ,n1167);
    or g1441(n1486 ,n1171 ,n1174);
    or g1442(n1485 ,n1179 ,n1166);
    or g1443(n1484 ,n1168 ,n1175);
    or g1444(n1483 ,n1160 ,n1172);
    or g1445(n1482 ,n1134 ,n1162);
    or g1446(n1481 ,n1159 ,n1156);
    or g1447(n1480 ,n1157 ,n1151);
    or g1448(n1479 ,n1155 ,n1153);
    or g1449(n1478 ,n959 ,n1325);
    or g1450(n1477 ,n1150 ,n1149);
    or g1451(n1476 ,n962 ,n1326);
    or g1452(n1475 ,n1146 ,n1145);
    or g1453(n1474 ,n1144 ,n1143);
    or g1454(n1473 ,n1142 ,n1138);
    nor g1455(n1472 ,n603 ,n1211);
    or g1456(n1471 ,n1137 ,n1136);
    or g1457(n1470 ,n1135 ,n1133);
    or g1458(n1469 ,n927 ,n1328);
    or g1459(n1468 ,n1141 ,n1208);
    or g1460(n1467 ,n1180 ,n1189);
    or g1461(n1466 ,n1169 ,n1209);
    or g1462(n1465 ,n1177 ,n1129);
    or g1463(n1464 ,n1214 ,n1128);
    nor g1464(n1463 ,n401 ,n1227);
    or g1465(n1462 ,n954 ,n1327);
    nor g1466(n1461 ,n203 ,n1140);
    or g1467(n1460 ,n1330 ,n1205);
    nor g1468(n1459 ,n6 ,n1212);
    or g1469(n1458 ,n1269 ,n1203);
    or g1470(n1457 ,n1307 ,n1193);
    or g1471(n1456 ,n1323 ,n1204);
    or g1472(n1455 ,n947 ,n1329);
    or g1473(n1454 ,n1301 ,n1201);
    or g1474(n1453 ,n1293 ,n1200);
    or g1475(n1452 ,n1343 ,n1199);
    or g1476(n1451 ,n1277 ,n1198);
    or g1477(n1450 ,n1306 ,n1197);
    or g1478(n1449 ,n1261 ,n1196);
    or g1479(n1448 ,n1253 ,n1195);
    or g1480(n1447 ,n1221 ,n1192);
    or g1481(n1446 ,n1245 ,n1194);
    or g1482(n1445 ,n1340 ,n1202);
    or g1483(n1444 ,n1303 ,n1191);
    or g1484(n1443 ,n934 ,n1335);
    or g1485(n1442 ,n926 ,n1334);
    or g1486(n1441 ,n929 ,n1333);
    or g1487(n1440 ,n1123 ,n1332);
    or g1488(n1439 ,n939 ,n1331);
    or g1489(n1438 ,n873 ,n1305);
    nor g1490(n1525 ,n203 ,n1230);
    or g1491(n1524 ,n229 ,n1213);
    nor g1492(n1522 ,n407 ,n1344);
    nor g1493(n1521 ,n669 ,n1229);
    nor g1494(n1518 ,n18[2] ,n1229);
    nor g1495(n1516 ,n675 ,n1344);
    not g1496(n1437 ,n1436);
    or g1497(n1435 ,n871 ,n1268);
    or g1498(n1434 ,n949 ,n1308);
    or g1499(n1433 ,n964 ,n1342);
    or g1500(n1432 ,n940 ,n1248);
    or g1501(n1431 ,n925 ,n1304);
    or g1502(n1430 ,n901 ,n1310);
    or g1503(n1429 ,n866 ,n1311);
    or g1504(n1428 ,n918 ,n1215);
    or g1505(n1427 ,n730 ,n1339);
    or g1506(n1426 ,n736 ,n1338);
    or g1507(n1425 ,n728 ,n1337);
    nor g1508(n1424 ,n666 ,n1228);
    or g1509(n1423 ,n922 ,n1216);
    nor g1510(n1422 ,n18[2] ,n1230);
    nor g1511(n1421 ,n18[1] ,n1207);
    or g1512(n1420 ,n879 ,n1316);
    or g1513(n1419 ,n909 ,n1300);
    or g1514(n1418 ,n951 ,n1299);
    or g1515(n1417 ,n894 ,n1298);
    or g1516(n1416 ,n892 ,n1297);
    or g1517(n1415 ,n890 ,n1296);
    or g1518(n1414 ,n906 ,n1295);
    or g1519(n1413 ,n880 ,n1294);
    or g1520(n1412 ,n899 ,n1292);
    or g1521(n1411 ,n887 ,n1291);
    or g1522(n1410 ,n963 ,n1290);
    or g1523(n1409 ,n885 ,n1289);
    or g1524(n1408 ,n908 ,n1288);
    or g1525(n1407 ,n898 ,n1314);
    or g1526(n1406 ,n928 ,n1287);
    or g1527(n1405 ,n893 ,n1286);
    or g1528(n1404 ,n923 ,n1284);
    or g1529(n1403 ,n886 ,n1283);
    or g1530(n1402 ,n881 ,n1282);
    or g1531(n1401 ,n883 ,n1281);
    or g1532(n1400 ,n903 ,n1280);
    or g1533(n1399 ,n889 ,n1218);
    or g1534(n1398 ,n904 ,n1279);
    or g1535(n1397 ,n849 ,n1278);
    or g1536(n1396 ,n865 ,n1276);
    or g1537(n1395 ,n874 ,n1275);
    or g1538(n1394 ,n930 ,n1274);
    or g1539(n1393 ,n875 ,n1273);
    or g1540(n1392 ,n958 ,n1272);
    or g1541(n1391 ,n936 ,n1271);
    or g1542(n1390 ,n955 ,n1270);
    or g1543(n1389 ,n952 ,n1309);
    or g1544(n1388 ,n900 ,n1267);
    or g1545(n1387 ,n946 ,n1266);
    or g1546(n1386 ,n919 ,n1265);
    or g1547(n1385 ,n985 ,n1264);
    or g1548(n1384 ,n912 ,n1263);
    or g1549(n1383 ,n852 ,n1262);
    or g1550(n1382 ,n867 ,n1260);
    or g1551(n1381 ,n861 ,n1259);
    or g1552(n1380 ,n864 ,n1258);
    or g1553(n1379 ,n857 ,n1257);
    or g1554(n1378 ,n916 ,n1256);
    or g1555(n1377 ,n882 ,n1255);
    or g1556(n1376 ,n920 ,n1254);
    or g1557(n1375 ,n917 ,n1252);
    or g1558(n1374 ,n937 ,n1251);
    or g1559(n1373 ,n935 ,n1250);
    or g1560(n1372 ,n944 ,n1249);
    or g1561(n1371 ,n948 ,n1247);
    or g1562(n1370 ,n957 ,n1246);
    or g1563(n1369 ,n984 ,n1244);
    or g1564(n1368 ,n858 ,n1243);
    or g1565(n1367 ,n897 ,n1242);
    or g1566(n1366 ,n986 ,n1241);
    or g1567(n1365 ,n956 ,n1240);
    or g1568(n1364 ,n941 ,n1239);
    or g1569(n1363 ,n913 ,n1238);
    or g1570(n1362 ,n950 ,n1236);
    or g1571(n1361 ,n856 ,n1235);
    or g1572(n1360 ,n878 ,n1234);
    or g1573(n1359 ,n905 ,n1233);
    or g1574(n1358 ,n933 ,n1232);
    or g1575(n1357 ,n855 ,n1285);
    or g1576(n1356 ,n961 ,n1336);
    or g1577(n1355 ,n921 ,n1319);
    or g1578(n1354 ,n896 ,n1237);
    or g1579(n1353 ,n938 ,n1341);
    or g1580(n1352 ,n850 ,n1225);
    or g1581(n1351 ,n860 ,n1223);
    or g1582(n1350 ,n851 ,n1222);
    or g1583(n1349 ,n960 ,n1224);
    or g1584(n1348 ,n872 ,n1220);
    or g1585(n1347 ,n877 ,n1219);
    or g1586(n1346 ,n884 ,n1217);
    or g1587(n1345 ,n891 ,n1302);
    nor g1588(n1436 ,n1148 ,n1206);
    nor g1589(n1343 ,n485 ,n979);
    nor g1590(n1342 ,n322 ,n968);
    nor g1591(n1341 ,n447 ,n968);
    nor g1592(n1340 ,n498 ,n968);
    nor g1593(n1339 ,n356 ,n981);
    nor g1594(n1338 ,n360 ,n981);
    nor g1595(n1337 ,n380 ,n981);
    nor g1596(n1336 ,n593 ,n974);
    nor g1597(n1335 ,n353 ,n971);
    nor g1598(n1334 ,n240 ,n971);
    nor g1599(n1333 ,n352 ,n971);
    nor g1600(n1332 ,n298 ,n971);
    nor g1601(n1331 ,n553 ,n971);
    nor g1602(n1330 ,n271 ,n967);
    nor g1603(n1329 ,n473 ,n967);
    nor g1604(n1328 ,n446 ,n967);
    nor g1605(n1327 ,n536 ,n967);
    nor g1606(n1326 ,n594 ,n967);
    nor g1607(n1325 ,n592 ,n967);
    nor g1608(n1324 ,n577 ,n967);
    nor g1609(n1323 ,n467 ,n970);
    nor g1610(n1322 ,n254 ,n970);
    nor g1611(n1321 ,n465 ,n970);
    nor g1612(n1320 ,n523 ,n970);
    nor g1613(n1319 ,n442 ,n970);
    nor g1614(n1318 ,n449 ,n970);
    nor g1615(n1317 ,n532 ,n970);
    nor g1616(n1316 ,n290 ,n970);
    nor g1617(n1315 ,n272 ,n973);
    nor g1618(n1314 ,n554 ,n973);
    nor g1619(n1313 ,n558 ,n973);
    nor g1620(n1312 ,n528 ,n973);
    nor g1621(n1311 ,n537 ,n973);
    nor g1622(n1310 ,n476 ,n973);
    nor g1623(n1309 ,n296 ,n973);
    nor g1624(n1308 ,n500 ,n967);
    nor g1625(n1307 ,n511 ,n974);
    nor g1626(n1306 ,n576 ,n977);
    nor g1627(n1305 ,n539 ,n971);
    nor g1628(n1304 ,n461 ,n971);
    nor g1629(n1303 ,n525 ,n971);
    nor g1630(n1302 ,n354 ,n972);
    nor g1631(n1301 ,n549 ,n966);
    nor g1632(n1300 ,n268 ,n966);
    nor g1633(n1299 ,n464 ,n966);
    nor g1634(n1298 ,n548 ,n966);
    nor g1635(n1297 ,n600 ,n966);
    nor g1636(n1296 ,n597 ,n966);
    nor g1637(n1295 ,n568 ,n966);
    nor g1638(n1294 ,n496 ,n966);
    nor g1639(n1293 ,n239 ,n980);
    nor g1640(n1292 ,n491 ,n980);
    nor g1641(n1291 ,n599 ,n980);
    nor g1642(n1290 ,n453 ,n980);
    nor g1643(n1289 ,n303 ,n980);
    nor g1644(n1288 ,n315 ,n980);
    nor g1645(n1287 ,n459 ,n980);
    nor g1646(n1286 ,n514 ,n980);
    nor g1647(n1285 ,n445 ,n974);
    nor g1648(n1284 ,n565 ,n979);
    nor g1649(n1283 ,n538 ,n979);
    nor g1650(n1282 ,n288 ,n979);
    nor g1651(n1281 ,n502 ,n979);
    nor g1652(n1280 ,n258 ,n979);
    nor g1653(n1279 ,n455 ,n979);
    nor g1654(n1278 ,n596 ,n979);
    nor g1655(n1277 ,n454 ,n978);
    nor g1656(n1276 ,n339 ,n978);
    nor g1657(n1275 ,n441 ,n978);
    nor g1658(n1274 ,n260 ,n978);
    nor g1659(n1273 ,n321 ,n978);
    nor g1660(n1272 ,n440 ,n978);
    nor g1661(n1271 ,n579 ,n978);
    nor g1662(n1270 ,n504 ,n978);
    nor g1663(n1269 ,n236 ,n973);
    nor g1664(n1268 ,n534 ,n977);
    nor g1665(n1267 ,n470 ,n977);
    nor g1666(n1266 ,n460 ,n977);
    nor g1667(n1265 ,n318 ,n977);
    nor g1668(n1264 ,n266 ,n977);
    nor g1669(n1263 ,n277 ,n977);
    nor g1670(n1262 ,n280 ,n977);
    nor g1671(n1261 ,n547 ,n976);
    nor g1672(n1260 ,n535 ,n976);
    nor g1673(n1259 ,n569 ,n976);
    nor g1674(n1258 ,n308 ,n976);
    nor g1675(n1257 ,n483 ,n976);
    nor g1676(n1256 ,n295 ,n976);
    nor g1677(n1255 ,n501 ,n976);
    nor g1678(n1254 ,n471 ,n976);
    nor g1679(n1253 ,n337 ,n969);
    nor g1680(n1252 ,n595 ,n969);
    nor g1681(n1251 ,n482 ,n969);
    nor g1682(n1250 ,n323 ,n969);
    nor g1683(n1249 ,n531 ,n969);
    nor g1684(n1248 ,n484 ,n969);
    nor g1685(n1247 ,n468 ,n969);
    nor g1686(n1246 ,n248 ,n969);
    nor g1687(n1245 ,n306 ,n975);
    nor g1688(n1244 ,n331 ,n975);
    nor g1689(n1243 ,n582 ,n975);
    nor g1690(n1242 ,n493 ,n975);
    nor g1691(n1241 ,n578 ,n975);
    nor g1692(n1240 ,n590 ,n975);
    nor g1693(n1239 ,n580 ,n975);
    nor g1694(n1238 ,n278 ,n975);
    nor g1695(n1237 ,n457 ,n968);
    nor g1696(n1236 ,n452 ,n974);
    nor g1697(n1235 ,n346 ,n974);
    nor g1698(n1234 ,n469 ,n974);
    nor g1699(n1233 ,n529 ,n974);
    nor g1700(n1232 ,n557 ,n974);
    or g1701(n1344 ,n223 ,n1124);
    not g1702(n1229 ,n1228);
    not g1703(n1227 ,n1226);
    nor g1704(n1225 ,n326 ,n968);
    nor g1705(n1224 ,n591 ,n968);
    nor g1706(n1223 ,n311 ,n968);
    nor g1707(n1222 ,n334 ,n968);
    nor g1708(n1221 ,n487 ,n972);
    nor g1709(n1220 ,n310 ,n972);
    nor g1710(n1219 ,n540 ,n972);
    nor g1711(n1218 ,n286 ,n972);
    nor g1712(n1217 ,n325 ,n972);
    nor g1713(n1216 ,n486 ,n972);
    nor g1714(n1215 ,n480 ,n972);
    or g1715(n1214 ,n1087 ,n1007);
    or g1716(n1213 ,n623 ,n1124);
    or g1717(n1212 ,n651 ,n1124);
    or g1718(n1211 ,n673 ,n1126);
    or g1719(n1210 ,n840 ,n994);
    or g1720(n1209 ,n1105 ,n1003);
    or g1721(n1208 ,n1012 ,n1011);
    nor g1722(n1207 ,n612 ,n1126);
    nor g1723(n1206 ,n401 ,n982);
    or g1724(n1205 ,n194 ,n943);
    or g1725(n1204 ,n194 ,n902);
    or g1726(n1203 ,n194 ,n876);
    or g1727(n1202 ,n200 ,n854);
    or g1728(n1201 ,n200 ,n895);
    or g1729(n1200 ,n195 ,n953);
    or g1730(n1199 ,n199 ,n910);
    or g1731(n1198 ,n202 ,n942);
    or g1732(n1197 ,n200 ,n870);
    or g1733(n1196 ,n200 ,n853);
    or g1734(n1195 ,n199 ,n914);
    or g1735(n1194 ,n195 ,n862);
    or g1736(n1193 ,n195 ,n932);
    or g1737(n1192 ,n195 ,n869);
    or g1738(n1191 ,n202 ,n924);
    or g1739(n1190 ,n1104 ,n1122);
    or g1740(n1189 ,n1005 ,n1108);
    or g1741(n1188 ,n783 ,n987);
    or g1742(n1187 ,n1117 ,n1081);
    or g1743(n1186 ,n1116 ,n1089);
    or g1744(n1185 ,n750 ,n1024);
    or g1745(n1184 ,n780 ,n988);
    or g1746(n1183 ,n781 ,n991);
    or g1747(n1182 ,n784 ,n989);
    or g1748(n1181 ,n1009 ,n1111);
    or g1749(n1180 ,n751 ,n1115);
    or g1750(n1179 ,n1085 ,n1079);
    or g1751(n1178 ,n779 ,n992);
    or g1752(n1177 ,n732 ,n1098);
    or g1753(n1176 ,n1004 ,n1006);
    or g1754(n1175 ,n1113 ,n1034);
    or g1755(n1174 ,n1099 ,n1101);
    or g1756(n1173 ,n777 ,n993);
    or g1757(n1172 ,n1084 ,n1082);
    or g1758(n1171 ,n1095 ,n1097);
    or g1759(n1170 ,n752 ,n1103);
    or g1760(n1169 ,n1107 ,n1102);
    or g1761(n1168 ,n1100 ,n1083);
    or g1762(n1167 ,n1121 ,n1076);
    or g1763(n1166 ,n1090 ,n1093);
    or g1764(n1165 ,n1072 ,n1086);
    or g1765(n1164 ,n778 ,n990);
    or g1766(n1163 ,n1013 ,n1118);
    or g1767(n1162 ,n1074 ,n1073);
    or g1768(n1161 ,n1071 ,n1070);
    or g1769(n1160 ,n1096 ,n1112);
    or g1770(n1159 ,n1065 ,n1064);
    or g1771(n1158 ,n998 ,n1066);
    or g1772(n1157 ,n734 ,n1061);
    or g1773(n1156 ,n1063 ,n1062);
    or g1774(n1155 ,n1060 ,n1059);
    or g1775(n1154 ,n1094 ,n1114);
    or g1776(n1153 ,n1058 ,n1056);
    or g1777(n1152 ,n1078 ,n1091);
    or g1778(n1151 ,n1057 ,n1054);
    or g1779(n1150 ,n735 ,n1053);
    or g1780(n1149 ,n1052 ,n1051);
    nor g1781(n1148 ,n18[1] ,n848);
    or g1782(n1147 ,n1049 ,n1048);
    or g1783(n1146 ,n1045 ,n1044);
    or g1784(n1145 ,n1042 ,n1041);
    or g1785(n1144 ,n1038 ,n1036);
    or g1786(n1143 ,n1120 ,n1035);
    or g1787(n1142 ,n1106 ,n1032);
    or g1788(n1141 ,n1015 ,n1014);
    nor g1789(n1140 ,n639 ,n844);
    or g1790(n1139 ,n620 ,n1125);
    or g1791(n1138 ,n1030 ,n1031);
    or g1792(n1137 ,n1029 ,n1039);
    or g1793(n1136 ,n1028 ,n1027);
    or g1794(n1135 ,n729 ,n1022);
    or g1795(n1134 ,n746 ,n1077);
    or g1796(n1133 ,n1025 ,n1023);
    or g1797(n1132 ,n1021 ,n1119);
    or g1798(n1131 ,n1050 ,n1047);
    or g1799(n1130 ,n1018 ,n1017);
    or g1800(n1129 ,n1020 ,n1068);
    or g1801(n1128 ,n1033 ,n1026);
    or g1802(n1127 ,n1016 ,n1037);
    or g1803(n1231 ,n690 ,n846);
    nor g1804(n1230 ,n1125 ,n847);
    nor g1805(n1228 ,n18[0] ,n1124);
    nor g1806(n1226 ,n407 ,n983);
    not g1807(n1126 ,n1125);
    nor g1808(n1123 ,n212 ,n827);
    nor g1809(n1122 ,n530 ,n834);
    nor g1810(n1121 ,n242 ,n833);
    nor g1811(n1120 ,n466 ,n802);
    nor g1812(n1119 ,n542 ,n837);
    nor g1813(n1118 ,n314 ,n804);
    nor g1814(n1117 ,n451 ,n805);
    nor g1815(n1116 ,n340 ,n835);
    nor g1816(n1115 ,n269 ,n832);
    nor g1817(n1114 ,n261 ,n800);
    nor g1818(n1113 ,n301 ,n799);
    nor g1819(n1112 ,n458 ,n803);
    nor g1820(n1111 ,n512 ,n801);
    nor g1821(n1110 ,n556 ,n836);
    nor g1822(n1109 ,n279 ,n836);
    nor g1823(n1108 ,n349 ,n834);
    nor g1824(n1107 ,n351 ,n839);
    nor g1825(n1106 ,n463 ,n839);
    nor g1826(n1105 ,n265 ,n799);
    nor g1827(n1104 ,n235 ,n833);
    nor g1828(n1103 ,n495 ,n832);
    nor g1829(n1102 ,n478 ,n801);
    nor g1830(n1101 ,n571 ,n804);
    nor g1831(n1100 ,n560 ,n839);
    nor g1832(n1099 ,n521 ,n799);
    nor g1833(n1098 ,n545 ,n832);
    nor g1834(n1097 ,n563 ,n801);
    nor g1835(n1096 ,n284 ,n805);
    nor g1836(n1095 ,n572 ,n839);
    nor g1837(n1094 ,n456 ,n802);
    nor g1838(n1093 ,n249 ,n800);
    nor g1839(n1092 ,n477 ,n836);
    nor g1840(n1091 ,n304 ,n837);
    nor g1841(n1090 ,n244 ,n802);
    nor g1842(n1089 ,n552 ,n837);
    nor g1843(n1088 ,n259 ,n838);
    nor g1844(n1087 ,n550 ,n805);
    nor g1845(n1086 ,n283 ,n837);
    nor g1846(n1085 ,n287 ,n805);
    nor g1847(n1084 ,n505 ,n802);
    nor g1848(n1083 ,n474 ,n801);
    nor g1849(n1082 ,n510 ,n800);
    nor g1850(n1081 ,n355 ,n803);
    nor g1851(n1080 ,n448 ,n838);
    nor g1852(n1079 ,n585 ,n803);
    nor g1853(n1078 ,n551 ,n835);
    nor g1854(n1077 ,n494 ,n832);
    nor g1855(n1076 ,n294 ,n834);
    nor g1856(n1075 ,n338 ,n838);
    nor g1857(n1074 ,n508 ,n833);
    nor g1858(n1073 ,n276 ,n834);
    nor g1859(n1072 ,n329 ,n835);
    nor g1860(n1071 ,n515 ,n835);
    nor g1861(n1070 ,n527 ,n837);
    nor g1862(n1069 ,n522 ,n836);
    nor g1863(n1068 ,n589 ,n834);
    nor g1864(n1067 ,n450 ,n836);
    nor g1865(n1066 ,n472 ,n838);
    nor g1866(n1065 ,n342 ,n839);
    nor g1867(n1064 ,n312 ,n801);
    nor g1868(n1063 ,n247 ,n799);
    nor g1869(n1062 ,n251 ,n804);
    nor g1870(n1061 ,n256 ,n832);
    nor g1871(n1060 ,n264 ,n805);
    nor g1872(n1059 ,n336 ,n803);
    nor g1873(n1058 ,n513 ,n802);
    nor g1874(n1057 ,n497 ,n833);
    nor g1875(n1056 ,n305 ,n800);
    nor g1876(n1055 ,n275 ,n838);
    nor g1877(n1054 ,n520 ,n834);
    nor g1878(n1053 ,n307 ,n832);
    nor g1879(n1052 ,n289 ,n833);
    nor g1880(n1051 ,n317 ,n834);
    nor g1881(n1050 ,n564 ,n835);
    nor g1882(n1049 ,n285 ,n835);
    nor g1883(n1048 ,n555 ,n837);
    nor g1884(n1047 ,n526 ,n837);
    nor g1885(n1046 ,n345 ,n836);
    nor g1886(n1045 ,n238 ,n839);
    nor g1887(n1044 ,n313 ,n801);
    nor g1888(n1043 ,n517 ,n836);
    nor g1889(n1042 ,n588 ,n799);
    nor g1890(n1041 ,n444 ,n804);
    nor g1891(n1040 ,n263 ,n838);
    nor g1892(n1039 ,n546 ,n803);
    nor g1893(n1038 ,n509 ,n805);
    nor g1894(n1037 ,n319 ,n804);
    nor g1895(n1036 ,n481 ,n803);
    nor g1896(n1035 ,n234 ,n800);
    nor g1897(n1034 ,n492 ,n804);
    nor g1898(n1033 ,n300 ,n802);
    nor g1899(n1032 ,n479 ,n801);
    nor g1900(n1031 ,n488 ,n804);
    nor g1901(n1030 ,n475 ,n799);
    nor g1902(n1029 ,n566 ,n805);
    nor g1903(n1028 ,n347 ,n802);
    nor g1904(n1027 ,n567 ,n800);
    nor g1905(n1026 ,n561 ,n800);
    nor g1906(n1025 ,n291 ,n833);
    nor g1907(n1024 ,n524 ,n832);
    nor g1908(n1023 ,n586 ,n834);
    nor g1909(n1022 ,n581 ,n832);
    nor g1910(n1021 ,n333 ,n835);
    nor g1911(n1020 ,n516 ,n833);
    nor g1912(n1019 ,n575 ,n836);
    nor g1913(n1018 ,n507 ,n839);
    nor g1914(n1017 ,n324 ,n801);
    nor g1915(n1016 ,n262 ,n799);
    nor g1916(n1015 ,n490 ,n805);
    nor g1917(n1014 ,n270 ,n803);
    nor g1918(n1013 ,n344 ,n799);
    nor g1919(n1012 ,n233 ,n802);
    nor g1920(n1011 ,n587 ,n800);
    nor g1921(n1010 ,n302 ,n838);
    nor g1922(n1009 ,n518 ,n839);
    nor g1923(n1008 ,n273 ,n838);
    nor g1924(n1007 ,n292 ,n803);
    nor g1925(n1006 ,n350 ,n837);
    nor g1926(n1005 ,n503 ,n833);
    nor g1927(n1004 ,n327 ,n835);
    nor g1928(n1003 ,n281 ,n804);
    nor g1929(n1002 ,n544 ,n825);
    nor g1930(n1001 ,n443 ,n825);
    nor g1931(n1000 ,n320 ,n825);
    nor g1932(n999 ,n559 ,n825);
    nor g1933(n998 ,n598 ,n825);
    nor g1934(n997 ,n237 ,n825);
    nor g1935(n996 ,n583 ,n825);
    nor g1936(n995 ,n584 ,n825);
    nor g1937(n994 ,n328 ,n806);
    nor g1938(n993 ,n499 ,n806);
    nor g1939(n992 ,n252 ,n806);
    nor g1940(n991 ,n533 ,n806);
    nor g1941(n990 ,n293 ,n806);
    nor g1942(n989 ,n348 ,n806);
    nor g1943(n988 ,n330 ,n806);
    nor g1944(n987 ,n245 ,n806);
    nor g1945(n986 ,n209 ,n811);
    nor g1946(n985 ,n212 ,n794);
    nor g1947(n984 ,n207 ,n811);
    nor g1948(n1125 ,n407 ,n831);
    or g1949(n1124 ,n421 ,n831);
    not g1950(n983 ,n982);
    nor g1951(n964 ,n208 ,n815);
    nor g1952(n963 ,n213 ,n819);
    nor g1953(n962 ,n209 ,n817);
    nor g1954(n961 ,n211 ,n823);
    nor g1955(n960 ,n209 ,n815);
    nor g1956(n959 ,n212 ,n817);
    nor g1957(n958 ,n212 ,n792);
    nor g1958(n957 ,n211 ,n829);
    nor g1959(n956 ,n212 ,n811);
    nor g1960(n955 ,n211 ,n792);
    nor g1961(n954 ,n214 ,n817);
    nor g1962(n953 ,n210 ,n819);
    nor g1963(n952 ,n211 ,n813);
    nor g1964(n951 ,n208 ,n788);
    nor g1965(n950 ,n207 ,n823);
    nor g1966(n949 ,n208 ,n817);
    nor g1967(n948 ,n214 ,n829);
    nor g1968(n947 ,n207 ,n817);
    nor g1969(n946 ,n213 ,n794);
    nor g1970(n945 ,n213 ,n796);
    nor g1971(n944 ,n209 ,n829);
    nor g1972(n943 ,n210 ,n817);
    nor g1973(n942 ,n210 ,n792);
    nor g1974(n941 ,n214 ,n811);
    nor g1975(n940 ,n212 ,n829);
    nor g1976(n939 ,n214 ,n827);
    nor g1977(n938 ,n207 ,n815);
    nor g1978(n937 ,n208 ,n829);
    nor g1979(n936 ,n214 ,n792);
    nor g1980(n935 ,n213 ,n829);
    nor g1981(n934 ,n207 ,n827);
    nor g1982(n933 ,n212 ,n823);
    nor g1983(n932 ,n210 ,n823);
    nor g1984(n931 ,n207 ,n796);
    nor g1985(n930 ,n213 ,n792);
    nor g1986(n929 ,n209 ,n827);
    nor g1987(n928 ,n214 ,n819);
    nor g1988(n927 ,n213 ,n817);
    nor g1989(n926 ,n213 ,n827);
    nor g1990(n925 ,n208 ,n827);
    nor g1991(n924 ,n210 ,n827);
    nor g1992(n923 ,n207 ,n790);
    nor g1993(n922 ,n214 ,n821);
    nor g1994(n921 ,n209 ,n796);
    nor g1995(n920 ,n211 ,n798);
    nor g1996(n919 ,n209 ,n794);
    nor g1997(n918 ,n211 ,n821);
    nor g1998(n917 ,n207 ,n829);
    nor g1999(n916 ,n212 ,n798);
    nor g2000(n915 ,n209 ,n813);
    nor g2001(n914 ,n210 ,n829);
    nor g2002(n913 ,n211 ,n811);
    nor g2003(n912 ,n214 ,n794);
    nor g2004(n911 ,n211 ,n817);
    nor g2005(n910 ,n210 ,n790);
    nor g2006(n909 ,n207 ,n788);
    nor g2007(n908 ,n212 ,n819);
    nor g2008(n907 ,n213 ,n813);
    nor g2009(n906 ,n214 ,n788);
    nor g2010(n905 ,n209 ,n823);
    nor g2011(n904 ,n214 ,n790);
    nor g2012(n903 ,n212 ,n790);
    nor g2013(n902 ,n210 ,n796);
    nor g2014(n901 ,n214 ,n813);
    nor g2015(n900 ,n208 ,n794);
    nor g2016(n899 ,n207 ,n819);
    nor g2017(n898 ,n208 ,n813);
    nor g2018(n897 ,n213 ,n811);
    nor g2019(n896 ,n212 ,n815);
    nor g2020(n895 ,n210 ,n788);
    nor g2021(n894 ,n213 ,n788);
    nor g2022(n893 ,n211 ,n819);
    nor g2023(n892 ,n209 ,n788);
    nor g2024(n891 ,n212 ,n821);
    nor g2025(n890 ,n212 ,n788);
    nor g2026(n889 ,n213 ,n821);
    nor g2027(n888 ,n207 ,n813);
    nor g2028(n887 ,n208 ,n819);
    nor g2029(n886 ,n208 ,n790);
    nor g2030(n885 ,n209 ,n819);
    nor g2031(n884 ,n209 ,n821);
    nor g2032(n883 ,n209 ,n790);
    nor g2033(n882 ,n214 ,n798);
    nor g2034(n881 ,n213 ,n790);
    nor g2035(n880 ,n211 ,n788);
    nor g2036(n879 ,n211 ,n796);
    nor g2037(n878 ,n213 ,n823);
    nor g2038(n877 ,n208 ,n821);
    nor g2039(n876 ,n210 ,n813);
    nor g2040(n875 ,n209 ,n792);
    nor g2041(n874 ,n208 ,n792);
    nor g2042(n873 ,n211 ,n827);
    nor g2043(n872 ,n207 ,n821);
    nor g2044(n871 ,n207 ,n794);
    nor g2045(n870 ,n210 ,n794);
    nor g2046(n869 ,n210 ,n821);
    nor g2047(n868 ,n214 ,n796);
    nor g2048(n867 ,n207 ,n798);
    nor g2049(n866 ,n212 ,n813);
    nor g2050(n865 ,n207 ,n792);
    nor g2051(n864 ,n213 ,n798);
    nor g2052(n863 ,n212 ,n796);
    nor g2053(n862 ,n210 ,n811);
    nor g2054(n861 ,n208 ,n798);
    nor g2055(n860 ,n214 ,n815);
    nor g2056(n859 ,n208 ,n796);
    nor g2057(n858 ,n208 ,n811);
    nor g2058(n857 ,n209 ,n798);
    nor g2059(n856 ,n208 ,n823);
    nor g2060(n855 ,n214 ,n823);
    nor g2061(n854 ,n210 ,n815);
    nor g2062(n853 ,n210 ,n798);
    nor g2063(n852 ,n211 ,n794);
    nor g2064(n851 ,n211 ,n815);
    nor g2065(n850 ,n213 ,n815);
    nor g2066(n849 ,n211 ,n790);
    nor g2067(n848 ,n203 ,n831);
    nor g2068(n847 ,n686 ,n831);
    nor g2069(n846 ,n671 ,n831);
    or g2070(n845 ,n716 ,n785);
    nor g2071(n844 ,n18[0] ,n831);
    or g2072(n843 ,n759 ,n808);
    or g2073(n842 ,n768 ,n807);
    or g2074(n841 ,n767 ,n809);
    or g2075(n840 ,n195 ,n782);
    nor g2076(n982 ,n18[2] ,n831);
    or g2077(n981 ,n713 ,n824);
    or g2078(n980 ,n194 ,n818);
    or g2079(n979 ,n201 ,n789);
    or g2080(n978 ,n201 ,n791);
    or g2081(n977 ,n199 ,n793);
    or g2082(n976 ,n201 ,n797);
    or g2083(n975 ,n202 ,n810);
    or g2084(n974 ,n200 ,n822);
    or g2085(n973 ,n200 ,n812);
    or g2086(n972 ,n199 ,n820);
    or g2087(n971 ,n202 ,n826);
    or g2088(n970 ,n194 ,n795);
    or g2089(n969 ,n194 ,n828);
    or g2090(n968 ,n200 ,n814);
    or g2091(n967 ,n200 ,n816);
    or g2092(n966 ,n195 ,n787);
    or g2093(n965 ,n745 ,n830);
    not g2094(n831 ,n830);
    not g2095(n829 ,n828);
    not g2096(n827 ,n826);
    not g2097(n825 ,n824);
    not g2098(n823 ,n822);
    not g2099(n821 ,n820);
    not g2100(n819 ,n818);
    not g2101(n817 ,n816);
    not g2102(n815 ,n814);
    not g2103(n813 ,n812);
    not g2104(n811 ,n810);
    nor g2105(n809 ,n358 ,n764);
    nor g2106(n808 ,n396 ,n764);
    nor g2107(n807 ,n388 ,n764);
    or g2108(n839 ,n647 ,n774);
    or g2109(n838 ,n645 ,n762);
    or g2110(n837 ,n642 ,n761);
    or g2111(n836 ,n642 ,n774);
    or g2112(n835 ,n642 ,n762);
    or g2113(n834 ,n645 ,n774);
    or g2114(n833 ,n645 ,n773);
    or g2115(n832 ,n647 ,n773);
    nor g2116(n830 ,n611 ,n757);
    nor g2117(n828 ,n681 ,n775);
    nor g2118(n826 ,n668 ,n776);
    nor g2119(n824 ,n642 ,n773);
    nor g2120(n822 ,n668 ,n766);
    nor g2121(n820 ,n668 ,n775);
    nor g2122(n818 ,n665 ,n765);
    nor g2123(n816 ,n682 ,n766);
    nor g2124(n814 ,n668 ,n765);
    nor g2125(n812 ,n682 ,n775);
    nor g2126(n810 ,n681 ,n776);
    not g2127(n798 ,n797);
    not g2128(n796 ,n795);
    not g2129(n794 ,n793);
    not g2130(n792 ,n791);
    not g2131(n790 ,n789);
    not g2132(n788 ,n787);
    nor g2133(n786 ,n197 ,n758);
    nor g2134(n785 ,n197 ,n755);
    nor g2135(n784 ,n214 ,n760);
    nor g2136(n783 ,n211 ,n760);
    nor g2137(n782 ,n210 ,n760);
    nor g2138(n781 ,n209 ,n760);
    nor g2139(n780 ,n208 ,n760);
    nor g2140(n779 ,n213 ,n760);
    nor g2141(n778 ,n212 ,n760);
    nor g2142(n777 ,n207 ,n760);
    nor g2143(n806 ,n739 ,n763);
    or g2144(n805 ,n616 ,n773);
    or g2145(n804 ,n647 ,n761);
    or g2146(n803 ,n616 ,n774);
    or g2147(n802 ,n616 ,n762);
    or g2148(n801 ,n645 ,n761);
    or g2149(n800 ,n616 ,n761);
    or g2150(n799 ,n647 ,n762);
    nor g2151(n797 ,n681 ,n765);
    nor g2152(n795 ,n682 ,n765);
    nor g2153(n793 ,n681 ,n766);
    nor g2154(n791 ,n665 ,n776);
    nor g2155(n789 ,n665 ,n775);
    nor g2156(n787 ,n665 ,n766);
    nor g2157(n772 ,n250 ,n738);
    nor g2158(n771 ,n241 ,n738);
    nor g2159(n770 ,n243 ,n738);
    nor g2160(n769 ,n274 ,n738);
    nor g2161(n768 ,n417 ,n740);
    nor g2162(n767 ,n215 ,n740);
    or g2163(n776 ,n408 ,n743);
    or g2164(n775 ,n408 ,n744);
    or g2165(n774 ,n413 ,n742);
    or g2166(n773 ,n413 ,n754);
    not g2167(n764 ,n763);
    nor g2168(n759 ,n408 ,n740);
    xnor g2169(n758 ,n726 ,n59[0]);
    or g2170(n757 ,n609 ,n731);
    or g2171(n756 ,n733 ,n741);
    or g2172(n755 ,n22[0] ,n745);
    or g2173(n766 ,n59[1] ,n744);
    or g2174(n765 ,n59[1] ,n743);
    nor g2175(n763 ,n683 ,n738);
    or g2176(n762 ,n39[1] ,n754);
    or g2177(n761 ,n39[1] ,n742);
    or g2178(n760 ,n684 ,n738);
    nor g2179(n753 ,n371 ,n713);
    nor g2180(n752 ,n570 ,n712);
    nor g2181(n751 ,n506 ,n712);
    nor g2182(n750 ,n255 ,n712);
    nor g2183(n749 ,n400 ,n713);
    nor g2184(n748 ,n359 ,n713);
    nor g2185(n747 ,n357 ,n713);
    nor g2186(n746 ,n282 ,n712);
    or g2187(n754 ,n422 ,n713);
    not g2188(n742 ,n741);
    not g2189(n740 ,n739);
    not g2190(n738 ,n737);
    nor g2191(n736 ,n416 ,n712);
    nor g2192(n735 ,n573 ,n712);
    nor g2193(n734 ,n309 ,n712);
    nor g2194(n733 ,n422 ,n712);
    nor g2195(n732 ,n341 ,n712);
    or g2196(n731 ,n676 ,n705);
    nor g2197(n730 ,n413 ,n712);
    nor g2198(n729 ,n297 ,n712);
    nor g2199(n728 ,n219 ,n712);
    nor g2200(n745 ,n688 ,n703);
    or g2201(n744 ,n59[0] ,n727);
    or g2202(n743 ,n419 ,n727);
    nor g2203(n741 ,n39[0] ,n713);
    nor g2204(n739 ,n196 ,n726);
    nor g2205(n737 ,n196 ,n727);
    not g2206(n727 ,n726);
    nor g2207(n725 ,n230 ,n695);
    nor g2208(n724 ,n232 ,n695);
    nor g2209(n723 ,n423 ,n695);
    nor g2210(n722 ,n225 ,n695);
    nor g2211(n721 ,n430 ,n695);
    nor g2212(n720 ,n439 ,n695);
    nor g2213(n719 ,n432 ,n695);
    nor g2214(n718 ,n224 ,n695);
    nor g2215(n717 ,n228 ,n695);
    nor g2216(n716 ,n420 ,n695);
    nor g2217(n715 ,n435 ,n695);
    nor g2218(n714 ,n425 ,n695);
    nor g2219(n726 ,n2561 ,n691);
    or g2220(n711 ,n635 ,n694);
    nor g2221(n710 ,n434 ,n695);
    nor g2222(n709 ,n431 ,n695);
    nor g2223(n708 ,n424 ,n695);
    nor g2224(n707 ,n222 ,n699);
    nor g2225(n706 ,n412 ,n696);
    or g2226(n705 ,n641 ,n693);
    nor g2227(n704 ,n426 ,n695);
    or g2228(n703 ,n659 ,n687);
    nor g2229(n702 ,n19[4] ,n699);
    nor g2230(n701 ,n20[4] ,n696);
    nor g2231(n700 ,n196 ,n689);
    or g2232(n713 ,n201 ,n698);
    or g2233(n712 ,n199 ,n697);
    not g2234(n698 ,n697);
    not g2235(n695 ,n694);
    or g2236(n693 ,n632 ,n678);
    or g2237(n699 ,n602 ,n664);
    nor g2238(n697 ,n343 ,n667);
    or g2239(n696 ,n607 ,n661);
    nor g2240(n694 ,n197 ,n663);
    or g2241(n691 ,n19[4] ,n667);
    or g2242(n690 ,n194 ,n666);
    nor g2243(n689 ,n625 ,n677);
    or g2244(n688 ,n628 ,n670);
    or g2245(n687 ,n625 ,n674);
    or g2246(n692 ,n672 ,n685);
    not g2247(n686 ,n685);
    not g2248(n684 ,n683);
    not g2249(n680 ,n679);
    or g2250(n678 ,n640 ,n606);
    nor g2251(n677 ,n429 ,n604);
    or g2252(n676 ,n601 ,n608);
    nor g2253(n685 ,n658 ,n638);
    nor g2254(n683 ,n637 ,n634);
    or g2255(n682 ,n215 ,n652);
    or g2256(n681 ,n215 ,n624);
    nor g2257(n679 ,n656 ,n643);
    not g2258(n675 ,n674);
    not g2259(n671 ,n670);
    not g2260(n667 ,n666);
    or g2261(n664 ,n19[1] ,n627);
    or g2262(n663 ,n401 ,n651);
    nor g2263(n662 ,n18[2] ,n610);
    or g2264(n661 ,n20[1] ,n626);
    nor g2265(n660 ,n401 ,n618);
    nor g2266(n659 ,n18[1] ,n651);
    nor g2267(n674 ,n18[0] ,n617);
    or g2268(n673 ,n194 ,n617);
    nor g2269(n672 ,n18[1] ,n630);
    nor g2270(n670 ,n401 ,n631);
    or g2271(n669 ,n4 ,n617);
    or g2272(n668 ,n59[2] ,n652);
    nor g2273(n666 ,n18[1] ,n619);
    or g2274(n665 ,n59[2] ,n624);
    or g2275(n641 ,n426 ,n439);
    or g2276(n640 ,n232 ,n424);
    nor g2277(n639 ,n407 ,n316);
    or g2278(n638 ,n216 ,n21[3]);
    or g2279(n637 ,n419 ,n408);
    nor g2280(n636 ,n429 ,n198);
    nor g2281(n635 ,n519 ,n198);
    or g2282(n634 ,n215 ,n417);
    or g2283(n633 ,n253 ,n4);
    or g2284(n632 ,n420 ,n22[1]);
    or g2285(n658 ,n409 ,n220);
    nor g2286(n657 ,n541 ,n196);
    or g2287(n656 ,n217 ,n418);
    nor g2288(n655 ,n332 ,n198);
    nor g2289(n654 ,n543 ,n197);
    or g2290(n653 ,n216 ,n21[0]);
    or g2291(n652 ,n417 ,n198);
    or g2292(n651 ,n407 ,n203);
    or g2293(n650 ,n411 ,n40[1]);
    or g2294(n649 ,n414 ,n40[2]);
    or g2295(n648 ,n415 ,n58[3]);
    or g2296(n647 ,n416 ,n39[3]);
    or g2297(n646 ,n218 ,n58[2]);
    or g2298(n645 ,n219 ,n39[2]);
    or g2299(n644 ,n414 ,n411);
    or g2300(n643 ,n415 ,n218);
    or g2301(n642 ,n416 ,n219);
    not g2302(n631 ,n630);
    not g2303(n629 ,n628);
    not g2304(n623 ,n622);
    not g2305(n619 ,n618);
    nor g2306(n613 ,n401 ,n197);
    nor g2307(n612 ,n203 ,n3);
    or g2308(n611 ,n22[12] ,n22[13]);
    nor g2309(n610 ,n18[0] ,n2);
    or g2310(n609 ,n22[14] ,n22[15]);
    or g2311(n608 ,n22[10] ,n22[11]);
    or g2312(n607 ,n20[2] ,n20[3]);
    or g2313(n606 ,n22[6] ,n22[7]);
    nor g2314(n605 ,n18[2] ,n2611);
    nor g2315(n604 ,n18[1] ,n18[2]);
    or g2316(n603 ,n4 ,n2612);
    or g2317(n602 ,n19[2] ,n19[3]);
    or g2318(n601 ,n22[8] ,n22[9]);
    nor g2319(n630 ,n203 ,n18[0]);
    nor g2320(n628 ,n401 ,n18[2]);
    or g2321(n627 ,n201 ,n19[0]);
    or g2322(n626 ,n194 ,n20[0]);
    nor g2323(n625 ,n18[2] ,n2563);
    or g2324(n624 ,n201 ,n59[3]);
    nor g2325(n622 ,n407 ,n197);
    or g2326(n621 ,n21[0] ,n21[2]);
    nor g2327(n620 ,n401 ,n203);
    nor g2328(n618 ,n18[0] ,n18[2]);
    or g2329(n617 ,n203 ,n18[1]);
    or g2330(n616 ,n39[2] ,n39[3]);
    or g2331(n615 ,n40[1] ,n40[2]);
    or g2332(n614 ,n58[2] ,n58[3]);
    not g2333(n600 ,n42[4]);
    not g2334(n599 ,n43[2]);
    not g2335(n598 ,n38[0]);
    not g2336(n597 ,n42[5]);
    not g2337(n596 ,n44[7]);
    not g2338(n595 ,n48[1]);
    not g2339(n594 ,n54[4]);
    not g2340(n593 ,n50[7]);
    not g2341(n592 ,n54[5]);
    not g2342(n591 ,n51[4]);
    not g2343(n590 ,n49[5]);
    not g2344(n589 ,n33[5]);
    not g2345(n588 ,n28[7]);
    not g2346(n587 ,n23[1]);
    not g2347(n586 ,n33[1]);
    not g2348(n585 ,n25[4]);
    not g2349(n584 ,n38[1]);
    not g2350(n583 ,n38[7]);
    not g2351(n582 ,n49[2]);
    not g2352(n581 ,n30[1]);
    not g2353(n580 ,n49[6]);
    not g2354(n579 ,n45[6]);
    not g2355(n578 ,n49[4]);
    not g2356(n577 ,n54[7]);
    not g2357(n576 ,n46[0]);
    not g2358(n575 ,n37[1]);
    not g2359(n574 ,n60[4]);
    not g2360(n573 ,n9[7]);
    not g2361(n572 ,n29[4]);
    not g2362(n571 ,n27[4]);
    not g2363(n570 ,n9[3]);
    not g2364(n569 ,n47[2]);
    not g2365(n568 ,n42[6]);
    not g2366(n567 ,n23[0]);
    not g2367(n566 ,n26[0]);
    not g2368(n565 ,n44[1]);
    not g2369(n564 ,n36[7]);
    not g2370(n563 ,n31[4]);
    not g2371(n562 ,n15);
    not g2372(n561 ,n23[2]);
    not g2373(n560 ,n29[5]);
    not g2374(n559 ,n38[2]);
    not g2375(n558 ,n56[3]);
    not g2376(n557 ,n50[5]);
    not g2377(n556 ,n37[2]);
    not g2378(n555 ,n35[0]);
    not g2379(n554 ,n56[2]);
    not g2380(n553 ,n53[6]);
    not g2381(n552 ,n35[3]);
    not g2382(n551 ,n36[5]);
    not g2383(n550 ,n26[2]);
    not g2384(n549 ,n42[0]);
    not g2385(n548 ,n42[3]);
    not g2386(n547 ,n47[0]);
    not g2387(n546 ,n25[0]);
    not g2388(n545 ,n30[5]);
    not g2389(n544 ,n38[4]);
    not g2390(n543 ,n17);
    not g2391(n542 ,n35[1]);
    not g2392(n541 ,n11[1]);
    not g2393(n540 ,n52[2]);
    not g2394(n539 ,n53[7]);
    not g2395(n538 ,n44[2]);
    not g2396(n537 ,n56[5]);
    not g2397(n536 ,n54[6]);
    not g2398(n535 ,n47[1]);
    not g2399(n534 ,n46[1]);
    not g2400(n533 ,n57[4]);
    not g2401(n532 ,n55[6]);
    not g2402(n531 ,n48[4]);
    not g2403(n530 ,n33[3]);
    not g2404(n529 ,n50[4]);
    not g2405(n528 ,n56[4]);
    not g2406(n527 ,n35[6]);
    not g2407(n526 ,n35[7]);
    not g2408(n525 ,n53[0]);
    not g2409(n524 ,n30[4]);
    not g2410(n523 ,n55[3]);
    not g2411(n522 ,n37[6]);
    not g2412(n521 ,n28[4]);
    not g2413(n520 ,n33[0]);
    not g2414(n519 ,n11[2]);
    not g2415(n518 ,n29[3]);
    not g2416(n517 ,n37[0]);
    not g2417(n516 ,n34[5]);
    not g2418(n515 ,n36[6]);
    not g2419(n514 ,n43[7]);
    not g2420(n513 ,n24[6]);
    not g2421(n512 ,n31[3]);
    not g2422(n511 ,n50[0]);
    not g2423(n510 ,n23[5]);
    not g2424(n509 ,n26[7]);
    not g2425(n508 ,n34[6]);
    not g2426(n507 ,n29[1]);
    not g2427(n506 ,n9[2]);
    not g2428(n505 ,n24[5]);
    not g2429(n504 ,n45[7]);
    not g2430(n503 ,n34[2]);
    not g2431(n502 ,n44[4]);
    not g2432(n501 ,n47[6]);
    not g2433(n500 ,n54[2]);
    not g2434(n499 ,n57[1]);
    not g2435(n498 ,n51[0]);
    not g2436(n497 ,n34[0]);
    not g2437(n496 ,n42[7]);
    not g2438(n495 ,n30[3]);
    not g2439(n494 ,n30[6]);
    not g2440(n493 ,n49[3]);
    not g2441(n492 ,n27[5]);
    not g2442(n491 ,n43[1]);
    not g2443(n490 ,n26[1]);
    not g2444(n489 ,n60[3]);
    not g2445(n488 ,n27[0]);
    not g2446(n487 ,n52[0]);
    not g2447(n486 ,n52[6]);
    not g2448(n485 ,n44[0]);
    not g2449(n484 ,n48[5]);
    not g2450(n483 ,n47[4]);
    not g2451(n482 ,n48[2]);
    not g2452(n481 ,n25[7]);
    not g2453(n480 ,n52[7]);
    not g2454(n479 ,n31[0]);
    not g2455(n478 ,n31[2]);
    not g2456(n477 ,n37[5]);
    not g2457(n476 ,n56[6]);
    not g2458(n475 ,n28[0]);
    not g2459(n474 ,n31[5]);
    not g2460(n473 ,n54[1]);
    not g2461(n472 ,n32[0]);
    not g2462(n471 ,n47[7]);
    not g2463(n470 ,n46[2]);
    not g2464(n469 ,n50[3]);
    not g2465(n468 ,n48[6]);
    not g2466(n467 ,n55[0]);
    not g2467(n466 ,n24[7]);
    not g2468(n465 ,n55[2]);
    not g2469(n464 ,n42[2]);
    not g2470(n463 ,n29[0]);
    not g2471(n462 ,n60[6]);
    not g2472(n461 ,n53[2]);
    not g2473(n460 ,n46[3]);
    not g2474(n459 ,n43[6]);
    not g2475(n458 ,n25[5]);
    not g2476(n457 ,n51[5]);
    not g2477(n456 ,n24[3]);
    not g2478(n455 ,n44[6]);
    not g2479(n454 ,n45[0]);
    not g2480(n453 ,n43[3]);
    not g2481(n452 ,n50[1]);
    not g2482(n451 ,n26[3]);
    not g2483(n450 ,n37[3]);
    not g2484(n449 ,n55[5]);
    not g2485(n448 ,n32[6]);
    not g2486(n447 ,n51[1]);
    not g2487(n446 ,n54[3]);
    not g2488(n445 ,n50[6]);
    not g2489(n444 ,n27[7]);
    not g2490(n443 ,n38[5]);
    not g2491(n442 ,n55[4]);
    not g2492(n441 ,n45[2]);
    not g2493(n440 ,n45[5]);
    not g2494(n439 ,n22[3]);
    not g2495(n438 ,n21[3]);
    not g2496(n437 ,n19[3]);
    not g2497(n436 ,n19[1]);
    not g2498(n435 ,n22[12]);
    not g2499(n434 ,n22[13]);
    not g2500(n433 ,n20[0]);
    not g2501(n432 ,n22[7]);
    not g2502(n431 ,n22[9]);
    not g2503(n430 ,n22[14]);
    not g2504(n429 ,n16);
    not g2505(n428 ,n19[0]);
    not g2506(n427 ,n19[2]);
    not g2507(n426 ,n22[2]);
    not g2508(n425 ,n22[8]);
    not g2509(n424 ,n22[5]);
    not g2510(n423 ,n22[11]);
    not g2511(n422 ,n39[0]);
    not g2512(n421 ,n14);
    not g2513(n420 ,n22[0]);
    not g2514(n419 ,n59[0]);
    not g2515(n418 ,n58[1]);
    not g2516(n417 ,n59[3]);
    not g2517(n416 ,n39[2]);
    not g2518(n415 ,n58[2]);
    not g2519(n414 ,n40[1]);
    not g2520(n413 ,n39[1]);
    not g2521(n412 ,n20[4]);
    not g2522(n411 ,n40[2]);
    not g2523(n410 ,n40[3]);
    not g2524(n409 ,n21[0]);
    not g2525(n408 ,n59[1]);
    not g2526(n407 ,n18[0]);
    not g2527(n406 ,n41[7]);
    not g2528(n405 ,n41[3]);
    not g2529(n404 ,n41[4]);
    not g2530(n403 ,n41[6]);
    not g2531(n402 ,n41[5]);
    not g2532(n401 ,n18[1]);
    not g2533(n400 ,n2608);
    not g2534(n399 ,n2590);
    not g2535(n398 ,n2589);
    not g2536(n397 ,n2592);
    not g2537(n396 ,n2564);
    not g2538(n395 ,n7[4]);
    not g2539(n394 ,n2582);
    not g2540(n393 ,n2570);
    not g2541(n392 ,n2578);
    not g2542(n391 ,n2584);
    not g2543(n390 ,n2574);
    not g2544(n389 ,n2586);
    not g2545(n388 ,n2566);
    not g2546(n387 ,n7[3]);
    not g2547(n386 ,n7[5]);
    not g2548(n385 ,n2577);
    not g2549(n384 ,n2595);
    not g2550(n383 ,n2588);
    not g2551(n382 ,n2596);
    not g2552(n381 ,n2575);
    not g2553(n380 ,n2569);
    not g2554(n379 ,n2573);
    not g2555(n378 ,n2579);
    not g2556(n377 ,n7[6]);
    not g2557(n376 ,n2594);
    not g2558(n375 ,n7[0]);
    not g2559(n374 ,n2585);
    not g2560(n373 ,n2581);
    not g2561(n372 ,n2593);
    not g2562(n371 ,n2607);
    not g2563(n370 ,n2572);
    not g2564(n369 ,n2580);
    not g2565(n368 ,n2587);
    not g2566(n367 ,n2571);
    not g2567(n366 ,n2583);
    not g2568(n365 ,n7[2]);
    not g2569(n364 ,n7[1]);
    not g2570(n363 ,n2591);
    not g2571(n362 ,n2576);
    not g2572(n361 ,n2597);
    not g2573(n360 ,n2568);
    not g2574(n359 ,n2609);
    not g2575(n358 ,n2565);
    not g2576(n357 ,n2610);
    not g2577(n356 ,n2567);
    not g2578(n355 ,n25[3]);
    not g2579(n354 ,n52[5]);
    not g2580(n353 ,n53[1]);
    not g2581(n352 ,n53[4]);
    not g2582(n351 ,n29[2]);
    not g2583(n350 ,n35[2]);
    not g2584(n349 ,n33[2]);
    not g2585(n348 ,n57[6]);
    not g2586(n347 ,n24[0]);
    not g2587(n346 ,n50[2]);
    not g2588(n345 ,n37[7]);
    not g2589(n344 ,n28[3]);
    not g2590(n343 ,n2611);
    not g2591(n342 ,n29[6]);
    not g2592(n341 ,n9[5]);
    not g2593(n340 ,n36[3]);
    not g2594(n339 ,n45[1]);
    not g2595(n338 ,n32[3]);
    not g2596(n337 ,n48[0]);
    not g2597(n336 ,n25[6]);
    not g2598(n335 ,n60[5]);
    not g2599(n334 ,n51[7]);
    not g2600(n333 ,n36[1]);
    not g2601(n332 ,n11[0]);
    not g2602(n331 ,n49[1]);
    not g2603(n330 ,n57[2]);
    not g2604(n329 ,n36[4]);
    not g2605(n328 ,n57[0]);
    not g2606(n327 ,n36[2]);
    not g2607(n326 ,n51[3]);
    not g2608(n325 ,n52[4]);
    not g2609(n324 ,n31[1]);
    not g2610(n323 ,n48[3]);
    not g2611(n322 ,n51[2]);
    not g2612(n321 ,n45[4]);
    not g2613(n320 ,n38[6]);
    not g2614(n319 ,n27[1]);
    not g2615(n318 ,n46[4]);
    not g2616(n317 ,n33[7]);
    not g2617(n316 ,n2);
    not g2618(n315 ,n43[5]);
    not g2619(n314 ,n27[3]);
    not g2620(n313 ,n31[7]);
    not g2621(n312 ,n31[6]);
    not g2622(n311 ,n51[6]);
    not g2623(n310 ,n52[1]);
    not g2624(n309 ,n9[0]);
    not g2625(n308 ,n47[3]);
    not g2626(n307 ,n30[7]);
    not g2627(n306 ,n49[0]);
    not g2628(n305 ,n23[6]);
    not g2629(n304 ,n35[5]);
    not g2630(n303 ,n43[4]);
    not g2631(n302 ,n32[2]);
    not g2632(n301 ,n28[5]);
    not g2633(n300 ,n24[2]);
    not g2634(n299 ,n60[1]);
    not g2635(n298 ,n53[5]);
    not g2636(n297 ,n9[1]);
    not g2637(n296 ,n56[7]);
    not g2638(n295 ,n47[5]);
    not g2639(n294 ,n33[4]);
    not g2640(n293 ,n57[5]);
    not g2641(n292 ,n25[2]);
    not g2642(n291 ,n34[1]);
    not g2643(n290 ,n55[7]);
    not g2644(n289 ,n34[7]);
    not g2645(n288 ,n44[3]);
    not g2646(n287 ,n26[4]);
    not g2647(n286 ,n52[3]);
    not g2648(n285 ,n36[0]);
    not g2649(n284 ,n26[5]);
    not g2650(n283 ,n35[4]);
    not g2651(n282 ,n9[6]);
    not g2652(n281 ,n27[2]);
    not g2653(n280 ,n46[7]);
    not g2654(n279 ,n37[4]);
    not g2655(n278 ,n49[7]);
    not g2656(n277 ,n46[6]);
    not g2657(n276 ,n33[6]);
    not g2658(n275 ,n32[7]);
    not g2659(n274 ,n2599);
    not g2660(n273 ,n32[5]);
    not g2661(n272 ,n56[1]);
    not g2662(n271 ,n54[0]);
    not g2663(n270 ,n25[1]);
    not g2664(n269 ,n30[2]);
    not g2665(n268 ,n42[1]);
    not g2666(n267 ,n60[2]);
    not g2667(n266 ,n46[5]);
    not g2668(n265 ,n28[2]);
    not g2669(n264 ,n26[6]);
    not g2670(n263 ,n32[1]);
    not g2671(n262 ,n28[1]);
    not g2672(n261 ,n23[3]);
    not g2673(n260 ,n45[3]);
    not g2674(n259 ,n32[4]);
    not g2675(n258 ,n44[5]);
    not g2676(n257 ,n60[7]);
    not g2677(n256 ,n30[0]);
    not g2678(n255 ,n9[4]);
    not g2679(n254 ,n55[1]);
    not g2680(n253 ,n2612);
    not g2681(n252 ,n57[3]);
    not g2682(n251 ,n27[6]);
    not g2683(n250 ,n2598);
    not g2684(n249 ,n23[4]);
    not g2685(n248 ,n48[7]);
    not g2686(n247 ,n28[6]);
    not g2687(n246 ,n60[0]);
    not g2688(n245 ,n57[7]);
    not g2689(n244 ,n24[4]);
    not g2690(n243 ,n2600);
    not g2691(n242 ,n34[4]);
    not g2692(n241 ,n2601);
    not g2693(n240 ,n53[3]);
    not g2694(n239 ,n43[0]);
    not g2695(n238 ,n29[7]);
    not g2696(n237 ,n38[3]);
    not g2697(n236 ,n56[0]);
    not g2698(n235 ,n34[3]);
    not g2699(n234 ,n23[7]);
    not g2700(n233 ,n24[1]);
    not g2701(n232 ,n22[4]);
    not g2702(n231 ,n20[1]);
    not g2703(n230 ,n22[10]);
    not g2704(n229 ,n6);
    not g2705(n228 ,n22[6]);
    not g2706(n227 ,n20[3]);
    not g2707(n226 ,n20[2]);
    not g2708(n225 ,n22[1]);
    not g2709(n224 ,n22[15]);
    not g2710(n223 ,n4);
    not g2711(n222 ,n19[4]);
    not g2712(n221 ,n40[0]);
    not g2713(n220 ,n21[1]);
    not g2714(n219 ,n39[3]);
    not g2715(n218 ,n58[3]);
    not g2716(n217 ,n58[0]);
    not g2717(n216 ,n21[2]);
    not g2718(n215 ,n59[2]);
    not g2719(n214 ,n8[6]);
    not g2720(n213 ,n8[3]);
    not g2721(n212 ,n8[5]);
    not g2722(n211 ,n8[7]);
    not g2723(n210 ,n8[0]);
    not g2724(n209 ,n8[4]);
    not g2725(n208 ,n8[2]);
    not g2726(n207 ,n8[1]);
    not g2727(n206 ,n41[2]);
    not g2728(n205 ,n41[0]);
    not g2729(n204 ,n41[1]);
    not g2730(n203 ,n18[2]);
    not g2731(n202 ,n1);
    not g2732(n201 ,n1);
    not g2733(n200 ,n1);
    not g2734(n199 ,n1);
    not g2735(n198 ,n1);
    not g2736(n197 ,n1);
    not g2737(n196 ,n1);
    not g2738(n195 ,n1);
    not g2739(n194 ,n1);
    or g2740(n193 ,n195 ,n965);
    or g2741(n192 ,n199 ,n965);
    or g2742(n191 ,n202 ,n965);
    or g2743(n190 ,n194 ,n965);
    or g2744(n189 ,n198 ,n965);
    or g2745(n188 ,n200 ,n965);
    or g2746(n187 ,n692 ,n1605);
    or g2747(n186 ,n221 ,n1624);
    xor g2748(n2597 ,n19[4] ,n70);
    xor g2749(n2596 ,n19[3] ,n68);
    nor g2750(n70 ,n19[3] ,n69);
    xor g2751(n2595 ,n19[2] ,n66);
    not g2752(n69 ,n68);
    nor g2753(n68 ,n19[2] ,n67);
    xnor g2754(n2594 ,n19[1] ,n19[0]);
    not g2755(n67 ,n66);
    nor g2756(n66 ,n19[1] ,n19[0]);
    xor g2757(n2610 ,n20[4] ,n65);
    xor g2758(n2609 ,n20[3] ,n63);
    nor g2759(n65 ,n20[3] ,n64);
    xor g2760(n2608 ,n20[2] ,n61);
    not g2761(n64 ,n63);
    nor g2762(n63 ,n20[2] ,n62);
    xnor g2763(n2607 ,n20[1] ,n20[0]);
    not g2764(n62 ,n61);
    nor g2765(n61 ,n20[1] ,n20[0]);
    or g2766(n2612 ,n72 ,n73);
    or g2767(n73 ,n19[3] ,n71);
    or g2768(n72 ,n19[2] ,n19[0]);
    or g2769(n71 ,n19[4] ,n19[1]);
    or g2770(n2611 ,n75 ,n76);
    or g2771(n76 ,n20[3] ,n74);
    or g2772(n75 ,n20[2] ,n20[0]);
    or g2773(n74 ,n20[4] ,n20[1]);
    xor g2774(n2601 ,n2606 ,n88);
    nor g2775(n2600 ,n87 ,n88);
    nor g2776(n88 ,n78 ,n86);
    nor g2777(n87 ,n2605 ,n85);
    nor g2778(n2598 ,n84 ,n85);
    not g2779(n86 ,n85);
    nor g2780(n85 ,n80 ,n83);
    nor g2781(n84 ,n2604 ,n82);
    nor g2782(n2599 ,n82 ,n81);
    not g2783(n83 ,n82);
    nor g2784(n82 ,n77 ,n79);
    nor g2785(n81 ,n2603 ,n2602);
    not g2786(n80 ,n2604);
    not g2787(n79 ,n2602);
    not g2788(n78 ,n2605);
    not g2789(n77 ,n2603);
    xor g2790(n2566 ,n59[3] ,n96);
    nor g2791(n2565 ,n95 ,n96);
    nor g2792(n96 ,n91 ,n94);
    nor g2793(n95 ,n59[2] ,n93);
    nor g2794(n2564 ,n93 ,n92);
    not g2795(n94 ,n93);
    nor g2796(n93 ,n89 ,n90);
    nor g2797(n92 ,n59[1] ,n59[0]);
    not g2798(n91 ,n59[2]);
    not g2799(n90 ,n59[0]);
    not g2800(n89 ,n59[1]);
    xor g2801(n2569 ,n39[3] ,n104);
    nor g2802(n2568 ,n103 ,n104);
    nor g2803(n104 ,n99 ,n102);
    nor g2804(n103 ,n39[2] ,n101);
    nor g2805(n2567 ,n101 ,n100);
    not g2806(n102 ,n101);
    nor g2807(n101 ,n97 ,n98);
    nor g2808(n100 ,n39[1] ,n39[0]);
    not g2809(n99 ,n39[2]);
    not g2810(n98 ,n39[0]);
    not g2811(n97 ,n39[1]);
    xor g2812(n2572 ,n58[3] ,n112);
    nor g2813(n2571 ,n111 ,n112);
    nor g2814(n112 ,n107 ,n110);
    nor g2815(n111 ,n58[2] ,n109);
    nor g2816(n2570 ,n109 ,n108);
    not g2817(n110 ,n109);
    nor g2818(n109 ,n105 ,n106);
    nor g2819(n108 ,n58[1] ,n58[0]);
    not g2820(n107 ,n58[2]);
    not g2821(n106 ,n58[0]);
    not g2822(n105 ,n58[1]);
    xor g2823(n2593 ,n22[15] ,n168);
    nor g2824(n2592 ,n167 ,n168);
    nor g2825(n168 ,n124 ,n166);
    nor g2826(n167 ,n22[14] ,n165);
    nor g2827(n2591 ,n164 ,n165);
    not g2828(n166 ,n165);
    nor g2829(n165 ,n114 ,n163);
    nor g2830(n164 ,n22[13] ,n162);
    nor g2831(n2590 ,n161 ,n162);
    not g2832(n163 ,n162);
    nor g2833(n162 ,n127 ,n160);
    nor g2834(n161 ,n22[12] ,n159);
    nor g2835(n2589 ,n158 ,n159);
    not g2836(n160 ,n159);
    nor g2837(n159 ,n123 ,n157);
    nor g2838(n158 ,n22[11] ,n156);
    nor g2839(n2588 ,n155 ,n156);
    not g2840(n157 ,n156);
    nor g2841(n156 ,n125 ,n154);
    nor g2842(n155 ,n22[10] ,n153);
    nor g2843(n2587 ,n152 ,n153);
    not g2844(n154 ,n153);
    nor g2845(n153 ,n122 ,n151);
    nor g2846(n152 ,n22[9] ,n150);
    nor g2847(n2586 ,n149 ,n150);
    not g2848(n151 ,n150);
    nor g2849(n150 ,n119 ,n148);
    nor g2850(n149 ,n22[8] ,n147);
    nor g2851(n2585 ,n146 ,n147);
    not g2852(n148 ,n147);
    nor g2853(n147 ,n120 ,n145);
    nor g2854(n146 ,n22[7] ,n144);
    nor g2855(n2584 ,n143 ,n144);
    not g2856(n145 ,n144);
    nor g2857(n144 ,n113 ,n142);
    nor g2858(n143 ,n22[6] ,n141);
    nor g2859(n2583 ,n140 ,n141);
    not g2860(n142 ,n141);
    nor g2861(n141 ,n118 ,n139);
    nor g2862(n140 ,n22[5] ,n138);
    nor g2863(n2582 ,n137 ,n138);
    not g2864(n139 ,n138);
    nor g2865(n138 ,n116 ,n136);
    nor g2866(n137 ,n22[4] ,n135);
    nor g2867(n2581 ,n134 ,n135);
    not g2868(n136 ,n135);
    nor g2869(n135 ,n115 ,n133);
    nor g2870(n134 ,n22[3] ,n132);
    nor g2871(n2580 ,n131 ,n132);
    not g2872(n133 ,n132);
    nor g2873(n132 ,n117 ,n130);
    nor g2874(n131 ,n22[2] ,n129);
    nor g2875(n2579 ,n129 ,n128);
    not g2876(n130 ,n129);
    nor g2877(n129 ,n121 ,n126);
    nor g2878(n128 ,n22[1] ,n22[0]);
    not g2879(n127 ,n22[12]);
    not g2880(n126 ,n22[0]);
    not g2881(n125 ,n22[10]);
    not g2882(n124 ,n22[14]);
    not g2883(n123 ,n22[11]);
    not g2884(n122 ,n22[9]);
    not g2885(n121 ,n22[1]);
    not g2886(n120 ,n22[7]);
    not g2887(n119 ,n22[8]);
    not g2888(n118 ,n22[5]);
    not g2889(n117 ,n22[2]);
    not g2890(n116 ,n22[4]);
    not g2891(n115 ,n22[3]);
    not g2892(n114 ,n22[13]);
    not g2893(n113 ,n22[6]);
    xor g2894(n2575 ,n21[3] ,n176);
    nor g2895(n2574 ,n175 ,n176);
    nor g2896(n176 ,n171 ,n174);
    nor g2897(n175 ,n21[2] ,n173);
    nor g2898(n2573 ,n173 ,n172);
    not g2899(n174 ,n173);
    nor g2900(n173 ,n169 ,n170);
    nor g2901(n172 ,n21[1] ,n21[0]);
    not g2902(n171 ,n21[2]);
    not g2903(n170 ,n21[0]);
    not g2904(n169 ,n21[1]);
    xor g2905(n2578 ,n40[3] ,n184);
    nor g2906(n2577 ,n183 ,n184);
    nor g2907(n184 ,n179 ,n182);
    nor g2908(n183 ,n40[2] ,n181);
    nor g2909(n2576 ,n181 ,n180);
    not g2910(n182 ,n181);
    nor g2911(n181 ,n177 ,n178);
    nor g2912(n180 ,n40[1] ,n40[0]);
    not g2913(n179 ,n40[2]);
    not g2914(n178 ,n40[0]);
    not g2915(n177 ,n40[1]);
    not g2916(n185 ,n1670);
endmodule
