module top(n0, n1, n2, n3, n4);
    input n0, n1;
    input [31:0] n2;
    input [3:0] n3;
    output [15:0] n4;
    wire n0, n1;
    wire [31:0] n2;
    wire [3:0] n3;
    wire [15:0] n4;
    wire [7:0] n5;
    wire [15:0] n6;
    wire [15:0] n7;
    wire [63:0] n8;
    wire [3:0] n9;
    wire [2:0] n10;
    wire [15:0] n11;
    wire [7:0] n12;
    wire [63:0] n13;
    wire [15:0] n14;
    wire n15, n16, n17, n18, n19, n20, n21, n22;
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    nor g0(n106 ,n11[11] ,n104);
    or g1(n18 ,n11[2] ,n11[1]);
    nor g2(n350 ,n88 ,n89);
    dff g3(.RN(n390), .SN(1'b1), .CK(n0), .D(n386), .Q(n13[12]));
    or g4(n209 ,n10[1] ,n205);
    dff g5(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n309), .Q(n6[7]));
    nor g6(n27 ,n15 ,n26);
    not g7(n39 ,n12[4]);
    not g8(n121 ,n370);
    dff g9(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n224), .Q(n11[6]));
    nor g10(n104 ,n73 ,n102);
    xor g11(n379 ,n8[37] ,n14[5]);
    dff g12(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n304), .Q(n6[10]));
    not g13(n125 ,n353);
    dff g14(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n200), .Q(n9[3]));
    nor g15(n355 ,n103 ,n104);
    not g16(n166 ,n12[3]);
    nor g17(n92 ,n61 ,n90);
    xor g18(n8[40] ,n2[8] ,n3[0]);
    xnor g19(n281 ,n278 ,n13[1]);
    not g20(n171 ,n9[1]);
    nor g21(n356 ,n106 ,n107);
    nor g22(n207 ,n177 ,n175);
    nor g23(n248 ,n146 ,n228);
    not g24(n155 ,n5[5]);
    nor g25(n324 ,n117 ,n320);
    xnor g26(n4[12] ,n338 ,n6[12]);
    nor g27(n316 ,n174 ,n297);
    nor g28(n224 ,n139 ,n186);
    dff g29(.RN(1'b1), .SN(n390), .CK(n0), .D(n14[10]), .Q(n14[11]));
    nor g30(n363 ,n59 ,n60);
    not g31(n135 ,n356);
    nor g32(n180 ,n152 ,n117);
    nor g33(n238 ,n157 ,n229);
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n195), .Q(n5[6]));
    nor g35(n179 ,n171 ,n117);
    nor g36(n225 ,n140 ,n186);
    dff g37(.RN(n390), .SN(1'b1), .CK(n0), .D(n387), .Q(n13[10]));
    nor g38(n368 ,n45 ,n44);
    not g39(n96 ,n95);
    nor g40(n277 ,n201 ,n276);
    nor g41(n351 ,n91 ,n92);
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n267), .Q(n12[7]));
    not g43(n108 ,n107);
    nor g44(n182 ,n123 ,n117);
    xor g45(n338 ,n337 ,n370);
    nor g46(n269 ,n117 ,n256);
    not g47(n170 ,n12[6]);
    xor g48(n383 ,n8[38] ,n14[6]);
    not g49(n87 ,n86);
    xor g50(n8[34] ,n2[2] ,n3[2]);
    xnor g51(n295 ,n278 ,n13[6]);
    nor g52(n266 ,n244 ,n262);
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n216), .Q(n11[11]));
    xor g54(n8[42] ,n2[10] ,n3[2]);
    not g55(n81 ,n80);
    dff g56(.RN(1'b1), .SN(n390), .CK(n0), .D(n14[2]), .Q(n14[3]));
    nor g57(n259 ,n236 ,n240);
    nor g58(n215 ,n138 ,n186);
    not g59(n55 ,n54);
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n226), .Q(n11[4]));
    nor g61(n274 ,n117 ,n253);
    not g62(n157 ,n12[4]);
    or g63(n24 ,n20 ,n23);
    not g64(n163 ,n5[1]);
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n198), .Q(n5[2]));
    dff g66(.RN(n390), .SN(1'b1), .CK(n0), .D(n14[7]), .Q(n14[8]));
    xnor g67(n4[9] ,n338 ,n6[9]);
    xnor g68(n380 ,n14[13] ,n14[15]);
    nor g69(n204 ,n151 ,n147);
    nor g70(n256 ,n249 ,n247);
    or g71(n232 ,n230 ,n231);
    not g72(n344 ,n369);
    dff g73(.RN(1'b1), .SN(n390), .CK(n0), .D(n14[11]), .Q(n14[12]));
    nor g74(n45 ,n41 ,n38);
    not g75(n296 ,n297);
    or g76(n361 ,n32 ,n36);
    xor g77(n8[38] ,n2[6] ,n3[2]);
    nor g78(n115 ,n11[14] ,n113);
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n193), .Q(n5[7]));
    dff g80(.RN(n390), .SN(1'b1), .CK(n0), .D(n371), .Q(n13[0]));
    not g81(n156 ,n7[5]);
    dff g82(.RN(n390), .SN(1'b1), .CK(n0), .D(n372), .Q(n13[4]));
    not g83(n153 ,n5[4]);
    xnor g84(n4[15] ,n338 ,n6[15]);
    nor g85(n311 ,n117 ,n294);
    not g86(n339 ,n5[3]);
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n220), .Q(n11[3]));
    nor g88(n195 ,n155 ,n117);
    nor g89(n317 ,n147 ,n296);
    nor g90(n217 ,n125 ,n186);
    nor g91(n91 ,n11[6] ,n89);
    nor g92(n353 ,n97 ,n98);
    nor g93(n193 ,n164 ,n117);
    xnor g94(n4[13] ,n338 ,n6[13]);
    nor g95(n359 ,n115 ,n116);
    nor g96(n255 ,n235 ,n233);
    not g97(n52 ,n51);
    not g98(n69 ,n11[1]);
    xnor g99(n337 ,n335 ,n332);
    not g100(n72 ,n11[14]);
    nor g101(n265 ,n10[2] ,n255);
    xor g102(n385 ,n8[45] ,n14[13]);
    not g103(n133 ,n349);
    nor g104(n112 ,n11[13] ,n110);
    xor g105(n376 ,n8[34] ,n14[2]);
    xnor g106(n332 ,n9[0] ,n10[0]);
    not g107(n90 ,n89);
    nor g108(n219 ,n137 ,n186);
    nor g109(n262 ,n10[2] ,n232);
    nor g110(n315 ,n250 ,n297);
    nor g111(n185 ,n156 ,n117);
    nor g112(n94 ,n11[7] ,n92);
    nor g113(n51 ,n40 ,n49);
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n301), .Q(n6[15]));
    nor g115(n243 ,n152 ,n228);
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n221), .Q(n11[2]));
    xnor g117(n4[1] ,n338 ,n6[1]);
    nor g118(n214 ,n142 ,n186);
    xor g119(n371 ,n8[32] ,n14[0]);
    or g120(n173 ,n7[5] ,n7[7]);
    nor g121(n213 ,n127 ,n186);
    nor g122(n247 ,n131 ,n228);
    or g123(n31 ,n12[2] ,n12[1]);
    nor g124(n230 ,n344 ,n188);
    not g125(n41 ,n12[1]);
    not g126(n99 ,n98);
    nor g127(n346 ,n77 ,n76);
    or g128(n201 ,n167 ,n123);
    nor g129(n48 ,n43 ,n46);
    dff g130(.RN(1'b1), .SN(n390), .CK(n0), .D(n14[6]), .Q(n14[7]));
    dff g131(.RN(n390), .SN(1'b1), .CK(n0), .D(n375), .Q(n13[3]));
    xor g132(n8[43] ,n2[11] ,n3[3]);
    not g133(n168 ,n9[2]);
    nor g134(n57 ,n42 ,n55);
    not g135(n154 ,n7[3]);
    xnor g136(n290 ,n278 ,n13[7]);
    xnor g137(n4[11] ,n338 ,n6[11]);
    nor g138(n323 ,n117 ,n322);
    not g139(n134 ,n367);
    not g140(n390 ,n1);
    dff g141(.RN(n390), .SN(1'b1), .CK(n0), .D(n376), .Q(n13[2]));
    nor g142(n191 ,n151 ,n117);
    not g143(n165 ,n12[5]);
    dff g144(.RN(n390), .SN(1'b1), .CK(n0), .D(n14[5]), .Q(n14[6]));
    or g145(n327 ,n339 ,n5[2]);
    xnor g146(n4[0] ,n338 ,n6[0]);
    nor g147(n77 ,n69 ,n74);
    not g148(n46 ,n45);
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n274), .Q(n12[0]));
    or g150(n334 ,n328 ,n333);
    xnor g151(n381 ,n14[10] ,n14[12]);
    not g152(n43 ,n12[2]);
    xnor g153(n4[6] ,n338 ,n6[6]);
    not g154(n123 ,n7[6]);
    nor g155(n216 ,n135 ,n186);
    not g156(n139 ,n351);
    nor g157(n242 ,n170 ,n229);
    not g158(n130 ,n362);
    not g159(n38 ,n12[0]);
    not g160(n158 ,n12[7]);
    nor g161(n319 ,n210 ,n297);
    xor g162(n8[44] ,n2[12] ,n3[0]);
    not g163(n63 ,n11[3]);
    not g164(n162 ,n12[1]);
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n303), .Q(n6[8]));
    xnor g166(n283 ,n278 ,n13[15]);
    nor g167(n197 ,n120 ,n117);
    or g168(n330 ,n343 ,n5[0]);
    nor g169(n107 ,n71 ,n105);
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n310), .Q(n6[6]));
    dff g171(.RN(n390), .SN(1'b1), .CK(n0), .D(n14[0]), .Q(n14[1]));
    xnor g172(n282 ,n278 ,n13[0]);
    nor g173(n244 ,n121 ,n228);
    not g174(n71 ,n11[11]);
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n272), .Q(n12[2]));
    xor g176(n374 ,n8[46] ,n14[14]);
    xor g177(n362 ,n12[7] ,n60);
    xor g178(n382 ,n8[39] ,n14[7]);
    or g179(n250 ,n10[2] ,n206);
    nor g180(n95 ,n68 ,n93);
    or g181(n210 ,n10[2] ,n188);
    xnor g182(n253 ,n229 ,n12[0]);
    nor g183(n223 ,n132 ,n186);
    nor g184(n59 ,n12[6] ,n57);
    dff g185(.RN(1'b1), .SN(n390), .CK(n0), .D(n389), .Q(n14[0]));
    not g186(n141 ,n359);
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n324), .Q(n10[2]));
    nor g188(n347 ,n79 ,n80);
    not g189(n161 ,n7[2]);
    dff g190(.RN(n390), .SN(1'b1), .CK(n0), .D(n14[12]), .Q(n14[13]));
    or g191(n22 ,n11[4] ,n21);
    nor g192(n246 ,n129 ,n228);
    not g193(n129 ,n363);
    not g194(n102 ,n101);
    or g195(n178 ,n161 ,n7[1]);
    not g196(n61 ,n11[6]);
    not g197(n132 ,n355);
    not g198(n146 ,n365);
    dff g199(.RN(1'b1), .SN(n390), .CK(n0), .D(n14[1]), .Q(n14[2]));
    dff g200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n197), .Q(n5[3]));
    xor g201(n375 ,n8[35] ,n14[3]);
    not g202(n136 ,n2[0]);
    nor g203(n348 ,n82 ,n83);
    nor g204(n325 ,n117 ,n321);
    xnor g205(n4[5] ,n338 ,n6[5]);
    nor g206(n97 ,n11[8] ,n95);
    or g207(n187 ,n10[0] ,n10[1]);
    xor g208(n8[46] ,n2[14] ,n3[2]);
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n223), .Q(n11[10]));
    not g210(n160 ,n7[1]);
    nor g211(n261 ,n237 ,n251);
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n312), .Q(n6[5]));
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n191), .Q(n7[1]));
    dff g214(.RN(n390), .SN(1'b1), .CK(n0), .D(n377), .Q(n13[11]));
    xnor g215(n292 ,n278 ,n13[5]);
    nor g216(n229 ,n148 ,n187);
    nor g217(n47 ,n12[2] ,n45);
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n189), .Q(n7[3]));
    nor g219(n54 ,n39 ,n52);
    not g220(n62 ,n11[13]);
    nor g221(n297 ,n266 ,n279);
    not g222(n145 ,n368);
    nor g223(n200 ,n168 ,n117);
    xor g224(n8[35] ,n2[3] ,n3[3]);
    dff g225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n271), .Q(n12[3]));
    nor g226(n237 ,n162 ,n229);
    xnor g227(n289 ,n278 ,n13[8]);
    nor g228(n231 ,n118 ,n187);
    or g229(n174 ,n10[0] ,n10[2]);
    xnor g230(n284 ,n278 ,n13[14]);
    dff g231(.RN(n390), .SN(1'b1), .CK(n0), .D(n379), .Q(n13[5]));
    nor g232(n354 ,n100 ,n101);
    nor g233(n199 ,n117 ,n119);
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n308), .Q(n6[13]));
    or g235(n16 ,n11[8] ,n11[7]);
    dff g236(.RN(1'b1), .SN(n390), .CK(n0), .D(n14[4]), .Q(n14[5]));
    nor g237(n184 ,n153 ,n117);
    nor g238(n116 ,n72 ,n114);
    nor g239(n176 ,n150 ,n10[0]);
    dff g240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n311), .Q(n6[3]));
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n179), .Q(n9[2]));
    not g242(n143 ,n346);
    not g243(n126 ,n347);
    not g244(n142 ,n358);
    nor g245(n239 ,n158 ,n229);
    nor g246(n226 ,n133 ,n186);
    nor g247(n190 ,n160 ,n117);
    nor g248(n82 ,n11[3] ,n80);
    dff g249(.RN(n390), .SN(1'b1), .CK(n0), .D(n374), .Q(n13[14]));
    dff g250(.RN(1'b1), .SN(n390), .CK(n0), .D(n14[9]), .Q(n14[10]));
    nor g251(n273 ,n117 ,n261);
    dff g252(.RN(n390), .SN(1'b1), .CK(n0), .D(n373), .Q(n13[15]));
    dff g253(.RN(1'b1), .SN(n390), .CK(n0), .D(n14[14]), .Q(n14[15]));
    nor g254(n305 ,n117 ,n287);
    or g255(n23 ,n11[5] ,n22);
    nor g256(n235 ,n149 ,n227);
    or g257(n35 ,n12[7] ,n34);
    not g258(n68 ,n11[7]);
    xor g259(n386 ,n8[44] ,n14[12]);
    not g260(n49 ,n48);
    not g261(n205 ,n204);
    nor g262(n300 ,n117 ,n282);
    not g263(n118 ,n3[0]);
    nor g264(n321 ,n314 ,n315);
    not g265(n37 ,n12[6]);
    or g266(n333 ,n330 ,n329);
    nor g267(n221 ,n126 ,n186);
    xor g268(n373 ,n8[47] ,n14[15]);
    not g269(n84 ,n83);
    or g270(n25 ,n11[0] ,n24);
    nor g271(n189 ,n161 ,n117);
    dff g272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n302), .Q(n6[14]));
    xnor g273(n4[3] ,n338 ,n6[3]);
    nor g274(n308 ,n117 ,n285);
    not g275(n164 ,n5[6]);
    dff g276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n300), .Q(n6[0]));
    nor g277(n192 ,n117 ,n136);
    nor g278(n357 ,n109 ,n110);
    dff g279(.RN(n390), .SN(1'b1), .CK(n0), .D(n14[3]), .Q(n14[4]));
    not g280(n122 ,n12[2]);
    nor g281(n183 ,n167 ,n117);
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n214), .Q(n11[13]));
    not g283(n117 ,n1);
    xnor g284(n4[4] ,n338 ,n6[4]);
    not g285(n228 ,n229);
    dff g286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n307), .Q(n6[9]));
    or g287(n202 ,n171 ,n168);
    not g288(n140 ,n354);
    nor g289(n198 ,n163 ,n117);
    xor g290(n360 ,n11[15] ,n116);
    not g291(n167 ,n7[4]);
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n313), .Q(n6[4]));
    nor g293(n307 ,n117 ,n291);
    not g294(n114 ,n113);
    or g295(n234 ,n7[3] ,n209);
    xor g296(n372 ,n8[36] ,n14[4]);
    xor g297(n8[33] ,n2[1] ,n3[1]);
    nor g298(n181 ,n117 ,n118);
    nor g299(n80 ,n65 ,n78);
    not g300(n152 ,n9[0]);
    xnor g301(n291 ,n278 ,n13[9]);
    not g302(n150 ,n11[0]);
    nor g303(n56 ,n12[5] ,n54);
    not g304(n93 ,n92);
    dff g305(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n305), .Q(n6[11]));
    dff g306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n219), .Q(n11[5]));
    nor g307(n257 ,n242 ,n246);
    nor g308(n60 ,n37 ,n58);
    not g309(n124 ,n348);
    xor g310(n377 ,n8[43] ,n14[11]);
    dff g311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n192), .Q(n7[0]));
    xor g312(n8[36] ,n2[4] ,n3[0]);
    not g313(n119 ,n13[0]);
    dff g314(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n306), .Q(n6[12]));
    nor g315(n175 ,n147 ,n370);
    nor g316(n320 ,n318 ,n319);
    nor g317(n177 ,n118 ,n10[0]);
    not g318(n151 ,n7[0]);
    not g319(n78 ,n77);
    nor g320(n98 ,n67 ,n96);
    xnor g321(n331 ,n11[0] ,n12[0]);
    dff g322(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n269), .Q(n12[5]));
    dff g323(.RN(n390), .SN(1'b1), .CK(n0), .D(n388), .Q(n13[9]));
    nor g324(n366 ,n50 ,n51);
    xnor g325(n4[7] ,n338 ,n6[7]);
    not g326(n75 ,n11[12]);
    nor g327(n349 ,n85 ,n86);
    or g328(n278 ,n243 ,n265);
    or g329(n369 ,n19 ,n29);
    nor g330(n304 ,n117 ,n280);
    dff g331(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n222), .Q(n11[1]));
    not g332(n30 ,n12[3]);
    nor g333(n26 ,n18 ,n25);
    not g334(n65 ,n11[2]);
    not g335(n105 ,n104);
    or g336(n336 ,n342 ,n334);
    nor g337(n218 ,n144 ,n186);
    xor g338(n8[41] ,n2[9] ,n3[1]);
    dff g339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n323), .Q(n10[0]));
    xnor g340(n294 ,n278 ,n13[3]);
    xor g341(n384 ,n8[40] ,n14[8]);
    nor g342(n89 ,n66 ,n87);
    dff g343(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n199), .Q(n5[0]));
    or g344(n186 ,n117 ,n118);
    dff g345(.RN(n390), .SN(1'b1), .CK(n0), .D(n378), .Q(n13[1]));
    not g346(n343 ,n361);
    not g347(n169 ,n5[0]);
    xnor g348(n335 ,n331 ,n7[0]);
    not g349(n111 ,n110);
    nor g350(n194 ,n169 ,n117);
    nor g351(n270 ,n117 ,n258);
    nor g352(n314 ,n149 ,n296);
    or g353(n36 ,n12[4] ,n35);
    nor g354(n236 ,n166 ,n229);
    not g355(n148 ,n10[2]);
    xnor g356(n285 ,n278 ,n13[13]);
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n273), .Q(n12[1]));
    not g358(n326 ,n9[0]);
    dff g359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n213), .Q(n11[15]));
    not g360(n128 ,n366);
    dff g361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n217), .Q(n11[8]));
    xnor g362(n280 ,n278 ,n13[10]);
    not g363(n66 ,n11[5]);
    xnor g364(n286 ,n278 ,n13[12]);
    or g365(n28 ,n11[15] ,n27);
    nor g366(n196 ,n159 ,n117);
    nor g367(n76 ,n11[1] ,n11[0]);
    nor g368(n358 ,n112 ,n113);
    dff g369(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n185), .Q(n7[6]));
    xor g370(n378 ,n8[33] ,n14[1]);
    dff g371(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n194), .Q(n5[1]));
    xor g372(n388 ,n8[41] ,n14[9]);
    xnor g373(n206 ,n149 ,n147);
    nor g374(n249 ,n165 ,n229);
    nor g375(n310 ,n117 ,n295);
    nor g376(n83 ,n63 ,n81);
    xor g377(n389 ,n380 ,n381);
    not g378(n64 ,n11[4]);
    nor g379(n271 ,n117 ,n259);
    or g380(n279 ,n275 ,n277);
    nor g381(n208 ,n11[0] ,n186);
    dff g382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n215), .Q(n11[12]));
    nor g383(n103 ,n11[10] ,n101);
    dff g384(.RN(1'b1), .SN(n390), .CK(n0), .D(n14[8]), .Q(n14[9]));
    xnor g385(n287 ,n278 ,n13[11]);
    dff g386(.RN(n390), .SN(1'b1), .CK(n0), .D(n385), .Q(n13[13]));
    nor g387(n88 ,n11[5] ,n86);
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n180), .Q(n9[1]));
    not g389(n172 ,n9[3]);
    nor g390(n254 ,n239 ,n245);
    nor g391(n352 ,n94 ,n95);
    xnor g392(n288 ,n278 ,n13[2]);
    not g393(n340 ,n5[7]);
    not g394(n149 ,n10[1]);
    dff g395(.RN(n390), .SN(1'b1), .CK(n0), .D(n384), .Q(n13[8]));
    xnor g396(n4[8] ,n338 ,n6[8]);
    nor g397(n113 ,n62 ,n111);
    nor g398(n268 ,n117 ,n257);
    or g399(n264 ,n172 ,n250);
    dff g400(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n325), .Q(n10[1]));
    not g401(n74 ,n11[0]);
    xor g402(n8[47] ,n2[15] ,n3[3]);
    nor g403(n53 ,n12[4] ,n51);
    nor g404(n364 ,n56 ,n57);
    nor g405(n267 ,n117 ,n254);
    dff g406(.RN(1'b1), .SN(n390), .CK(n0), .D(n14[13]), .Q(n14[14]));
    or g407(n328 ,n340 ,n5[6]);
    nor g408(n367 ,n47 ,n48);
    nor g409(n245 ,n130 ,n228);
    nor g410(n212 ,n141 ,n186);
    dff g411(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n183), .Q(n7[5]));
    nor g412(n101 ,n70 ,n99);
    xnor g413(n293 ,n278 ,n13[4]);
    nor g414(n306 ,n117 ,n286);
    dff g415(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n225), .Q(n11[9]));
    nor g416(n241 ,n122 ,n229);
    not g417(n120 ,n5[2]);
    nor g418(n309 ,n117 ,n290);
    or g419(n19 ,n11[14] ,n11[13]);
    nor g420(n86 ,n64 ,n84);
    xor g421(n8[39] ,n2[7] ,n3[3]);
    nor g422(n258 ,n238 ,n248);
    nor g423(n44 ,n12[1] ,n12[0]);
    nor g424(n227 ,n204 ,n176);
    nor g425(n272 ,n117 ,n260);
    dff g426(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n212), .Q(n11[14]));
    nor g427(n50 ,n12[3] ,n48);
    xor g428(n387 ,n8[42] ,n14[10]);
    dff g429(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n181), .Q(n9[0]));
    nor g430(n233 ,n10[1] ,n207);
    not g431(n147 ,n10[0]);
    not g432(n42 ,n12[5]);
    xor g433(n8[32] ,n2[0] ,n3[0]);
    or g434(n21 ,n17 ,n16);
    dff g435(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n298), .Q(n6[2]));
    or g436(n211 ,n345 ,n202);
    nor g437(n313 ,n117 ,n293);
    nor g438(n34 ,n30 ,n33);
    nor g439(n318 ,n148 ,n296);
    xor g440(n8[37] ,n2[5] ,n3[1]);
    not g441(n70 ,n11[9]);
    not g442(n127 ,n360);
    nor g443(n100 ,n11[9] ,n98);
    not g444(n73 ,n11[10]);
    dff g445(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n196), .Q(n5[4]));
    dff g446(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n270), .Q(n12[4]));
    not g447(n144 ,n352);
    nor g448(n312 ,n117 ,n292);
    nor g449(n252 ,n134 ,n228);
    nor g450(n79 ,n11[2] ,n77);
    nor g451(n301 ,n117 ,n283);
    not g452(n15 ,n11[11]);
    nor g453(n260 ,n241 ,n252);
    not g454(n341 ,n5[5]);
    nor g455(n222 ,n143 ,n186);
    nor g456(n251 ,n145 ,n228);
    nor g457(n110 ,n75 ,n108);
    dff g458(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n208), .Q(n11[0]));
    xnor g459(n4[14] ,n338 ,n6[14]);
    nor g460(n299 ,n117 ,n281);
    nor g461(n302 ,n117 ,n284);
    or g462(n276 ,n178 ,n263);
    nor g463(n220 ,n124 ,n186);
    nor g464(n203 ,n154 ,n117);
    not g465(n342 ,n5[1]);
    nor g466(n109 ,n11[12] ,n107);
    nor g467(n240 ,n128 ,n228);
    nor g468(n85 ,n11[4] ,n83);
    dff g469(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n184), .Q(n5[5]));
    nor g470(n33 ,n12[0] ,n31);
    dff g471(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n299), .Q(n6[1]));
    or g472(n345 ,n326 ,n10[0]);
    not g473(n137 ,n350);
    or g474(n17 ,n11[10] ,n11[9]);
    not g475(n67 ,n11[8]);
    not g476(n40 ,n12[3]);
    not g477(n138 ,n357);
    dff g478(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n218), .Q(n11[7]));
    dff g479(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n182), .Q(n7[7]));
    dff g480(.RN(n390), .SN(1'b1), .CK(n0), .D(n383), .Q(n13[6]));
    or g481(n263 ,n173 ,n234);
    dff g482(.RN(n390), .SN(1'b1), .CK(n0), .D(n382), .Q(n13[7]));
    or g483(n188 ,n147 ,n149);
    or g484(n32 ,n12[6] ,n12[5]);
    xnor g485(n4[2] ,n338 ,n6[2]);
    nor g486(n365 ,n53 ,n54);
    xor g487(n8[45] ,n2[13] ,n3[1]);
    not g488(n159 ,n5[3]);
    dff g489(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n268), .Q(n12[6]));
    not g490(n131 ,n364);
    not g491(n58 ,n57);
    or g492(n370 ,n327 ,n336);
    or g493(n29 ,n11[12] ,n28);
    dff g494(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n203), .Q(n7[4]));
    nor g495(n322 ,n317 ,n316);
    or g496(n20 ,n11[6] ,n11[3]);
    nor g497(n275 ,n211 ,n264);
    or g498(n329 ,n341 ,n5[4]);
    xnor g499(n4[10] ,n338 ,n6[10]);
    dff g500(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n190), .Q(n7[2]));
    nor g501(n298 ,n117 ,n288);
    nor g502(n303 ,n117 ,n289);
endmodule
