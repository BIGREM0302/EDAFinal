module top(n0, n1, n4, n6, n5, n2, n11, n12, n13, n14, n17, n15, n16, n3, n7, n8, n9, n10);
    input n0, n1, n2, n3;
    input [7:0] n4;
    input [3:0] n5;
    output [7:0] n6, n7, n8, n9, n10;
    output n11, n12, n13, n14, n15, n16;
    output [3:0] n17;
    wire n0, n1, n2, n3;
    wire [7:0] n4;
    wire [3:0] n5;
    wire [7:0] n6, n7, n8, n9, n10;
    wire n11, n12, n13, n14, n15, n16;
    wire [3:0] n17;
    wire [3:0] n18;
    wire [3:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [7:0] n22;
    wire [7:0] n23;
    wire [7:0] n24;
    wire [7:0] n25;
    wire [7:0] n26;
    wire [7:0] n27;
    wire [7:0] n28;
    wire [7:0] n29;
    wire [7:0] n30;
    wire [7:0] n31;
    wire [7:0] n32;
    wire [7:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [4:0] n36;
    wire [3:0] n37;
    wire [3:0] n38;
    wire [7:0] n39;
    wire [2:0] n40;
    wire [7:0] n41;
    wire [7:0] n42;
    wire [7:0] n43;
    wire [7:0] n44;
    wire [7:0] n45;
    wire [7:0] n46;
    wire [7:0] n47;
    wire [7:0] n48;
    wire [7:0] n49;
    wire [7:0] n50;
    wire [7:0] n51;
    wire [7:0] n52;
    wire [7:0] n53;
    wire [7:0] n54;
    wire [7:0] n55;
    wire [7:0] n56;
    wire [4:0] n57;
    wire [3:0] n58;
    wire [3:0] n59;
    wire [7:0] n60;
    wire n61, n62, n63, n64, n65, n66, n67, n68;
    wire n69, n70, n71, n72, n73, n74, n75, n76;
    wire n77, n78, n79, n80, n81, n82, n83, n84;
    wire n85, n86, n87, n88, n89, n90, n91, n92;
    wire n93, n94, n95, n96, n97, n98, n99, n100;
    wire n101, n102, n103, n104, n105, n106, n107, n108;
    wire n109, n110, n111, n112, n113, n114, n115, n116;
    wire n117, n118, n119, n120, n121, n122, n123, n124;
    wire n125, n126, n127, n128, n129, n130, n131, n132;
    wire n133, n134, n135, n136, n137, n138, n139, n140;
    wire n141, n142, n143, n144, n145, n146, n147, n148;
    wire n149, n150, n151, n152, n153, n154, n155, n156;
    wire n157, n158, n159, n160, n161, n162, n163, n164;
    wire n165, n166, n167, n168, n169, n170, n171, n172;
    wire n173, n174, n175, n176, n177, n178, n179, n180;
    wire n181, n182, n183, n184, n185, n186, n187, n188;
    wire n189, n190, n191, n192, n193, n194, n195, n196;
    wire n197, n198, n199, n200, n201, n202, n203, n204;
    wire n205, n206, n207, n208, n209, n210, n211, n212;
    wire n213, n214, n215, n216, n217, n218, n219, n220;
    wire n221, n222, n223, n224, n225, n226, n227, n228;
    wire n229, n230, n231, n232, n233, n234, n235, n236;
    wire n237, n238, n239, n240, n241, n242, n243, n244;
    wire n245, n246, n247, n248, n249, n250, n251, n252;
    wire n253, n254, n255, n256, n257, n258, n259, n260;
    wire n261, n262, n263, n264, n265, n266, n267, n268;
    wire n269, n270, n271, n272, n273, n274, n275, n276;
    wire n277, n278, n279, n280, n281, n282, n283, n284;
    wire n285, n286, n287, n288, n289, n290, n291, n292;
    wire n293, n294, n295, n296, n297, n298, n299, n300;
    wire n301, n302, n303, n304, n305, n306, n307, n308;
    wire n309, n310, n311, n312, n313, n314, n315, n316;
    wire n317, n318, n319, n320, n321, n322, n323, n324;
    wire n325, n326, n327, n328, n329, n330, n331, n332;
    wire n333, n334, n335, n336, n337, n338, n339, n340;
    wire n341, n342, n343, n344, n345, n346, n347, n348;
    wire n349, n350, n351, n352, n353, n354, n355, n356;
    wire n357, n358, n359, n360, n361, n362, n363, n364;
    wire n365, n366, n367, n368, n369, n370, n371, n372;
    wire n373, n374, n375, n376, n377, n378, n379, n380;
    wire n381, n382, n383, n384, n385, n386, n387, n388;
    wire n389, n390, n391, n392, n393, n394, n395, n396;
    wire n397, n398, n399, n400, n401, n402, n403, n404;
    wire n405, n406, n407, n408, n409, n410, n411, n412;
    wire n413, n414, n415, n416, n417, n418, n419, n420;
    wire n421, n422, n423, n424, n425, n426, n427, n428;
    wire n429, n430, n431, n432, n433, n434, n435, n436;
    wire n437, n438, n439, n440, n441, n442, n443, n444;
    wire n445, n446, n447, n448, n449, n450, n451, n452;
    wire n453, n454, n455, n456, n457, n458, n459, n460;
    wire n461, n462, n463, n464, n465, n466, n467, n468;
    wire n469, n470, n471, n472, n473, n474, n475, n476;
    wire n477, n478, n479, n480, n481, n482, n483, n484;
    wire n485, n486, n487, n488, n489, n490, n491, n492;
    wire n493, n494, n495, n496, n497, n498, n499, n500;
    wire n501, n502, n503, n504, n505, n506, n507, n508;
    wire n509, n510, n511, n512, n513, n514, n515, n516;
    wire n517, n518, n519, n520, n521, n522, n523, n524;
    wire n525, n526, n527, n528, n529, n530, n531, n532;
    wire n533, n534, n535, n536, n537, n538, n539, n540;
    wire n541, n542, n543, n544, n545, n546, n547, n548;
    wire n549, n550, n551, n552, n553, n554, n555, n556;
    wire n557, n558, n559, n560, n561, n562, n563, n564;
    wire n565, n566, n567, n568, n569, n570, n571, n572;
    wire n573, n574, n575, n576, n577, n578, n579, n580;
    wire n581, n582, n583, n584, n585, n586, n587, n588;
    wire n589, n590, n591, n592, n593, n594, n595, n596;
    wire n597, n598, n599, n600, n601, n602, n603, n604;
    wire n605, n606, n607, n608, n609, n610, n611, n612;
    wire n613, n614, n615, n616, n617, n618, n619, n620;
    wire n621, n622, n623, n624, n625, n626, n627, n628;
    wire n629, n630, n631, n632, n633, n634, n635, n636;
    wire n637, n638, n639, n640, n641, n642, n643, n644;
    wire n645, n646, n647, n648, n649, n650, n651, n652;
    wire n653, n654, n655, n656, n657, n658, n659, n660;
    wire n661, n662, n663, n664, n665, n666, n667, n668;
    wire n669, n670, n671, n672, n673, n674, n675, n676;
    wire n677, n678, n679, n680, n681, n682, n683, n684;
    wire n685, n686, n687, n688, n689, n690, n691, n692;
    wire n693, n694, n695, n696, n697, n698, n699, n700;
    wire n701, n702, n703, n704, n705, n706, n707, n708;
    wire n709, n710, n711, n712, n713, n714, n715, n716;
    wire n717, n718, n719, n720, n721, n722, n723, n724;
    wire n725, n726, n727, n728, n729, n730, n731, n732;
    wire n733, n734, n735, n736, n737, n738, n739, n740;
    wire n741, n742, n743, n744, n745, n746, n747, n748;
    wire n749, n750, n751, n752, n753, n754, n755, n756;
    wire n757, n758, n759, n760, n761, n762, n763, n764;
    wire n765, n766, n767, n768, n769, n770, n771, n772;
    wire n773, n774, n775, n776, n777, n778, n779, n780;
    wire n781, n782, n783, n784, n785, n786, n787, n788;
    wire n789, n790, n791, n792, n793, n794, n795, n796;
    wire n797, n798, n799, n800, n801, n802, n803, n804;
    wire n805, n806, n807, n808, n809, n810, n811, n812;
    wire n813, n814, n815, n816, n817, n818, n819, n820;
    wire n821, n822, n823, n824, n825, n826, n827, n828;
    wire n829, n830, n831, n832, n833, n834, n835, n836;
    wire n837, n838, n839, n840, n841, n842, n843, n844;
    wire n845, n846, n847, n848, n849, n850, n851, n852;
    wire n853, n854, n855, n856, n857, n858, n859, n860;
    wire n861, n862, n863, n864, n865, n866, n867, n868;
    wire n869, n870, n871, n872, n873, n874, n875, n876;
    wire n877, n878, n879, n880, n881, n882, n883, n884;
    wire n885, n886, n887, n888, n889, n890, n891, n892;
    wire n893, n894, n895, n896, n897, n898, n899, n900;
    wire n901, n902, n903, n904, n905, n906, n907, n908;
    wire n909, n910, n911, n912, n913, n914, n915, n916;
    wire n917, n918, n919, n920, n921, n922, n923, n924;
    wire n925, n926, n927, n928, n929, n930, n931, n932;
    wire n933, n934, n935, n936, n937, n938, n939, n940;
    wire n941, n942, n943, n944, n945, n946, n947, n948;
    wire n949, n950, n951, n952, n953, n954, n955, n956;
    wire n957, n958, n959, n960, n961, n962, n963, n964;
    wire n965, n966, n967, n968, n969, n970, n971, n972;
    wire n973, n974, n975, n976, n977, n978, n979, n980;
    wire n981, n982, n983, n984, n985, n986, n987, n988;
    wire n989, n990, n991, n992, n993, n994, n995, n996;
    wire n997, n998, n999, n1000, n1001, n1002, n1003, n1004;
    wire n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012;
    wire n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
    wire n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
    wire n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
    wire n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044;
    wire n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052;
    wire n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060;
    wire n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068;
    wire n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076;
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084;
    wire n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092;
    wire n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100;
    wire n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108;
    wire n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116;
    wire n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124;
    wire n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132;
    wire n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140;
    wire n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148;
    wire n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156;
    wire n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164;
    wire n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172;
    wire n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180;
    wire n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188;
    wire n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196;
    wire n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204;
    wire n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
    wire n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220;
    wire n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228;
    wire n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236;
    wire n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244;
    wire n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252;
    wire n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260;
    wire n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268;
    wire n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276;
    wire n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284;
    wire n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292;
    wire n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300;
    wire n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308;
    wire n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;
    wire n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;
    wire n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332;
    wire n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340;
    wire n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348;
    wire n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356;
    wire n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364;
    wire n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372;
    wire n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380;
    wire n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388;
    wire n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396;
    wire n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404;
    wire n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412;
    wire n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420;
    wire n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428;
    wire n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436;
    wire n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444;
    wire n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452;
    wire n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460;
    wire n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468;
    wire n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476;
    wire n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484;
    wire n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492;
    wire n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500;
    wire n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508;
    wire n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516;
    wire n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524;
    wire n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532;
    wire n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540;
    wire n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548;
    wire n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556;
    wire n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564;
    wire n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572;
    wire n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580;
    wire n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588;
    wire n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596;
    wire n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604;
    wire n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612;
    wire n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620;
    wire n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628;
    wire n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636;
    wire n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644;
    wire n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652;
    wire n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660;
    wire n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668;
    wire n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676;
    wire n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684;
    wire n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692;
    wire n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700;
    wire n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708;
    wire n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716;
    wire n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724;
    wire n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732;
    wire n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740;
    wire n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748;
    wire n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756;
    wire n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764;
    wire n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772;
    wire n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780;
    wire n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788;
    wire n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796;
    wire n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804;
    wire n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812;
    wire n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820;
    wire n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828;
    wire n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836;
    wire n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844;
    wire n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852;
    wire n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860;
    wire n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868;
    wire n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876;
    wire n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884;
    wire n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892;
    wire n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900;
    wire n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908;
    wire n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916;
    wire n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924;
    wire n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932;
    wire n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940;
    wire n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948;
    wire n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956;
    wire n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964;
    wire n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972;
    wire n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980;
    wire n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988;
    wire n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996;
    wire n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004;
    wire n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012;
    wire n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020;
    wire n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028;
    wire n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036;
    wire n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044;
    wire n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052;
    wire n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060;
    wire n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068;
    wire n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076;
    wire n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084;
    wire n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092;
    wire n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100;
    wire n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108;
    wire n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116;
    wire n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124;
    wire n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132;
    wire n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140;
    wire n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148;
    wire n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156;
    wire n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164;
    wire n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172;
    wire n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180;
    wire n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188;
    wire n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196;
    wire n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204;
    wire n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212;
    wire n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220;
    wire n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228;
    wire n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236;
    wire n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244;
    wire n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252;
    wire n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260;
    wire n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268;
    wire n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276;
    wire n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284;
    wire n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292;
    wire n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300;
    wire n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308;
    wire n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316;
    wire n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324;
    wire n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332;
    wire n2333;
    buf g0(n10[0], 1'b0);
    buf g1(n10[1], 1'b0);
    buf g2(n10[2], 1'b0);
    buf g3(n10[3], n7[1]);
    buf g4(n10[4], n7[7]);
    buf g5(n10[5], n7[7]);
    buf g6(n9[0], 1'b0);
    buf g7(n9[1], 1'b0);
    buf g8(n9[2], 1'b0);
    buf g9(n9[3], 1'b0);
    buf g10(n9[4], 1'b0);
    buf g11(n9[5], 1'b0);
    buf g12(n9[6], 1'b0);
    buf g13(n9[7], 1'b0);
    buf g14(n8[0], 1'b0);
    buf g15(n8[2], 1'b0);
    buf g16(n8[3], 1'b0);
    buf g17(n8[4], 1'b0);
    buf g18(n8[5], 1'b0);
    buf g19(n8[6], 1'b0);
    buf g20(n8[7], 1'b0);
    buf g21(n7[0], 1'b0);
    buf g22(n7[6], n7[7]);
    buf g23(n14, n13);
    not g24(n2299 ,n2333);
    not g25(n2298 ,n2332);
    not g26(n2297 ,n2316);
    not g27(n2296 ,n3);
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1270), .Q(n18[0]));
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1240), .Q(n18[1]));
    dff g30(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1398), .Q(n18[2]));
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1406), .Q(n18[3]));
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n606), .Q(n19[0]));
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n665), .Q(n19[1]));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n911), .Q(n17[0]));
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n912), .Q(n17[1]));
    dff g36(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n913), .Q(n17[2]));
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n914), .Q(n17[3]));
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n546), .Q(n7[1]));
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n530), .Q(n7[7]));
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n525), .Q(n10[6]));
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n519), .Q(n10[7]));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1879), .Q(n8[1]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n917), .Q(n16));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n576), .Q(n13));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2272), .Q(n6[0]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2276), .Q(n6[1]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2269), .Q(n6[2]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2267), .Q(n6[3]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2266), .Q(n6[4]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2265), .Q(n6[5]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2279), .Q(n6[6]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2274), .Q(n6[7]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2168), .Q(n12));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2184), .Q(n20[0]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2133), .Q(n20[1]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2132), .Q(n20[2]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2131), .Q(n20[3]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2130), .Q(n20[4]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2129), .Q(n20[5]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2128), .Q(n20[6]));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2127), .Q(n20[7]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2183), .Q(n21[0]));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2126), .Q(n21[1]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2125), .Q(n21[2]));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2124), .Q(n21[3]));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2123), .Q(n21[4]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2122), .Q(n21[5]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2121), .Q(n21[6]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2120), .Q(n21[7]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2181), .Q(n22[0]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2119), .Q(n22[1]));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2118), .Q(n22[2]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2117), .Q(n22[3]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2116), .Q(n22[4]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2115), .Q(n22[5]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2114), .Q(n22[6]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2113), .Q(n22[7]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2180), .Q(n23[0]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2112), .Q(n23[1]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2111), .Q(n23[2]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2110), .Q(n23[3]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2109), .Q(n23[4]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2108), .Q(n23[5]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2107), .Q(n23[6]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2106), .Q(n23[7]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2179), .Q(n24[0]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2105), .Q(n24[1]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2104), .Q(n24[2]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2103), .Q(n24[3]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2102), .Q(n24[4]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2101), .Q(n24[5]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2100), .Q(n24[6]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2099), .Q(n24[7]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2177), .Q(n25[0]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2098), .Q(n25[1]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2097), .Q(n25[2]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2096), .Q(n25[3]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2095), .Q(n25[4]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2094), .Q(n25[5]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2093), .Q(n25[6]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2092), .Q(n25[7]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2176), .Q(n26[0]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2091), .Q(n26[1]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2090), .Q(n26[2]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2089), .Q(n26[3]));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2088), .Q(n26[4]));
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2087), .Q(n26[5]));
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2086), .Q(n26[6]));
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2085), .Q(n26[7]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2175), .Q(n27[0]));
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2084), .Q(n27[1]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2083), .Q(n27[2]));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2082), .Q(n27[3]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2081), .Q(n27[4]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2080), .Q(n27[5]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2079), .Q(n27[6]));
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2078), .Q(n27[7]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2174), .Q(n28[0]));
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2077), .Q(n28[1]));
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2076), .Q(n28[2]));
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2075), .Q(n28[3]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2074), .Q(n28[4]));
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2073), .Q(n28[5]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2072), .Q(n28[6]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2071), .Q(n28[7]));
    dff g126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2171), .Q(n29[0]));
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2070), .Q(n29[1]));
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2069), .Q(n29[2]));
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2068), .Q(n29[3]));
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2067), .Q(n29[4]));
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2066), .Q(n29[5]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2065), .Q(n29[6]));
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2064), .Q(n29[7]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2169), .Q(n30[0]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2063), .Q(n30[1]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2140), .Q(n30[2]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2167), .Q(n30[3]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2166), .Q(n30[4]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2165), .Q(n30[5]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2164), .Q(n30[6]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2163), .Q(n30[7]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2196), .Q(n31[0]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2162), .Q(n31[1]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2161), .Q(n31[2]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2160), .Q(n31[3]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2159), .Q(n31[4]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2158), .Q(n31[5]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2157), .Q(n31[6]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2156), .Q(n31[7]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2195), .Q(n32[0]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2155), .Q(n32[1]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2154), .Q(n32[2]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2153), .Q(n32[3]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2152), .Q(n32[4]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2151), .Q(n32[5]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2150), .Q(n32[6]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2149), .Q(n32[7]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2193), .Q(n33[0]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2148), .Q(n33[1]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2147), .Q(n33[2]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2146), .Q(n33[3]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2145), .Q(n33[4]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2143), .Q(n33[5]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2144), .Q(n33[6]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2142), .Q(n33[7]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2192), .Q(n34[0]));
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2141), .Q(n34[1]));
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2208), .Q(n34[2]));
    dff g169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2209), .Q(n34[3]));
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2210), .Q(n34[4]));
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2211), .Q(n34[5]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2212), .Q(n34[6]));
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2213), .Q(n34[7]));
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2190), .Q(n35[0]));
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2062), .Q(n35[1]));
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2139), .Q(n35[2]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2138), .Q(n35[3]));
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2137), .Q(n35[4]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2136), .Q(n35[5]));
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2135), .Q(n35[6]));
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2134), .Q(n35[7]));
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1878), .Q(n36[0]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2188), .Q(n36[1]));
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2187), .Q(n36[2]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2186), .Q(n36[3]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2185), .Q(n36[4]));
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n684), .Q(n37[0]));
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1658), .Q(n37[1]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1659), .Q(n37[2]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1660), .Q(n37[3]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1894), .Q(n38[0]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2216), .Q(n38[1]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2215), .Q(n38[2]));
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2214), .Q(n38[3]));
    dff g195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1379), .Q(n39[0]));
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1378), .Q(n39[1]));
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1377), .Q(n39[2]));
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1375), .Q(n39[3]));
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1374), .Q(n39[4]));
    dff g200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1373), .Q(n39[5]));
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1372), .Q(n39[6]));
    dff g202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n685), .Q(n15));
    dff g203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1661), .Q(n40[0]));
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1663), .Q(n40[1]));
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n661), .Q(n7[2]));
    dff g206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n666), .Q(n7[3]));
    dff g207(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n619), .Q(n7[4]));
    dff g208(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n621), .Q(n7[5]));
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n916), .Q(n11));
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1685), .Q(n41[0]));
    dff g211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1366), .Q(n41[1]));
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1365), .Q(n41[2]));
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1363), .Q(n41[3]));
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1361), .Q(n41[4]));
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1360), .Q(n41[5]));
    dff g216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1359), .Q(n41[6]));
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1357), .Q(n41[7]));
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1684), .Q(n42[0]));
    dff g219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1355), .Q(n42[1]));
    dff g220(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1354), .Q(n42[2]));
    dff g221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1353), .Q(n42[3]));
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1352), .Q(n42[4]));
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1351), .Q(n42[5]));
    dff g224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1350), .Q(n42[6]));
    dff g225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1349), .Q(n42[7]));
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1683), .Q(n43[0]));
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1346), .Q(n43[1]));
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1345), .Q(n43[2]));
    dff g229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1343), .Q(n43[3]));
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1341), .Q(n43[4]));
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1340), .Q(n43[5]));
    dff g232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1339), .Q(n43[6]));
    dff g233(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1338), .Q(n43[7]));
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1682), .Q(n44[0]));
    dff g235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1337), .Q(n44[1]));
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1336), .Q(n44[2]));
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1335), .Q(n44[3]));
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1334), .Q(n44[4]));
    dff g239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1333), .Q(n44[5]));
    dff g240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1332), .Q(n44[6]));
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1331), .Q(n44[7]));
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1681), .Q(n45[0]));
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1328), .Q(n45[1]));
    dff g244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1327), .Q(n45[2]));
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1326), .Q(n45[3]));
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1324), .Q(n45[4]));
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1323), .Q(n45[5]));
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1322), .Q(n45[6]));
    dff g249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1321), .Q(n45[7]));
    dff g250(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1680), .Q(n46[0]));
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1318), .Q(n46[1]));
    dff g252(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1317), .Q(n46[2]));
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1315), .Q(n46[3]));
    dff g254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1314), .Q(n46[4]));
    dff g255(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1312), .Q(n46[5]));
    dff g256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1311), .Q(n46[6]));
    dff g257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1310), .Q(n46[7]));
    dff g258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1679), .Q(n47[0]));
    dff g259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1309), .Q(n47[1]));
    dff g260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1307), .Q(n47[2]));
    dff g261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1306), .Q(n47[3]));
    dff g262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1305), .Q(n47[4]));
    dff g263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1304), .Q(n47[5]));
    dff g264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1302), .Q(n47[6]));
    dff g265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1301), .Q(n47[7]));
    dff g266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1678), .Q(n48[0]));
    dff g267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1298), .Q(n48[1]));
    dff g268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1297), .Q(n48[2]));
    dff g269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1296), .Q(n48[3]));
    dff g270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1295), .Q(n48[4]));
    dff g271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1293), .Q(n48[5]));
    dff g272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1291), .Q(n48[6]));
    dff g273(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1290), .Q(n48[7]));
    dff g274(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1677), .Q(n49[0]));
    dff g275(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1288), .Q(n49[1]));
    dff g276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1286), .Q(n49[2]));
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1284), .Q(n49[3]));
    dff g278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1282), .Q(n49[4]));
    dff g279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1281), .Q(n49[5]));
    dff g280(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1280), .Q(n49[6]));
    dff g281(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1278), .Q(n49[7]));
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1676), .Q(n50[0]));
    dff g283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1276), .Q(n50[1]));
    dff g284(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1275), .Q(n50[2]));
    dff g285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1274), .Q(n50[3]));
    dff g286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1273), .Q(n50[4]));
    dff g287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1272), .Q(n50[5]));
    dff g288(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1271), .Q(n50[6]));
    dff g289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1269), .Q(n50[7]));
    dff g290(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1675), .Q(n51[0]));
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1267), .Q(n51[1]));
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1266), .Q(n51[2]));
    dff g293(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1264), .Q(n51[3]));
    dff g294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1362), .Q(n51[4]));
    dff g295(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1262), .Q(n51[5]));
    dff g296(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1261), .Q(n51[6]));
    dff g297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1397), .Q(n51[7]));
    dff g298(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1674), .Q(n52[0]));
    dff g299(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1257), .Q(n52[1]));
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1255), .Q(n52[2]));
    dff g301(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1371), .Q(n52[3]));
    dff g302(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1253), .Q(n52[4]));
    dff g303(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1283), .Q(n52[5]));
    dff g304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1252), .Q(n52[6]));
    dff g305(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1251), .Q(n52[7]));
    dff g306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1673), .Q(n53[0]));
    dff g307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1249), .Q(n53[1]));
    dff g308(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1248), .Q(n53[2]));
    dff g309(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1247), .Q(n53[3]));
    dff g310(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1246), .Q(n53[4]));
    dff g311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1245), .Q(n53[5]));
    dff g312(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1244), .Q(n53[6]));
    dff g313(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1242), .Q(n53[7]));
    dff g314(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1672), .Q(n54[0]));
    dff g315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1263), .Q(n54[1]));
    dff g316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1300), .Q(n54[2]));
    dff g317(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1239), .Q(n54[3]));
    dff g318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1238), .Q(n54[4]));
    dff g319(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1237), .Q(n54[5]));
    dff g320(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1316), .Q(n54[6]));
    dff g321(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1319), .Q(n54[7]));
    dff g322(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1671), .Q(n55[0]));
    dff g323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1234), .Q(n55[1]));
    dff g324(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1232), .Q(n55[2]));
    dff g325(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1368), .Q(n55[3]));
    dff g326(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1387), .Q(n55[4]));
    dff g327(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1230), .Q(n55[5]));
    dff g328(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1390), .Q(n55[6]));
    dff g329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1229), .Q(n55[7]));
    dff g330(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1688), .Q(n56[0]));
    dff g331(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1381), .Q(n56[1]));
    dff g332(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1409), .Q(n56[2]));
    dff g333(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1407), .Q(n56[3]));
    dff g334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1405), .Q(n56[4]));
    dff g335(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1404), .Q(n56[5]));
    dff g336(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1402), .Q(n56[6]));
    dff g337(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1401), .Q(n56[7]));
    dff g338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1400), .Q(n57[0]));
    dff g339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1414), .Q(n57[1]));
    dff g340(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1418), .Q(n57[2]));
    dff g341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1417), .Q(n57[3]));
    dff g342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1415), .Q(n57[4]));
    dff g343(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n921), .Q(n58[0]));
    dff g344(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1882), .Q(n58[1]));
    dff g345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1881), .Q(n58[2]));
    dff g346(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1880), .Q(n58[3]));
    dff g347(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1396), .Q(n59[0]));
    dff g348(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1653), .Q(n59[1]));
    dff g349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1652), .Q(n59[2]));
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1651), .Q(n59[3]));
    dff g351(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2284), .Q(n60[0]));
    dff g352(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2294), .Q(n60[1]));
    dff g353(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2295), .Q(n60[2]));
    dff g354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2293), .Q(n60[3]));
    dff g355(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2290), .Q(n60[4]));
    dff g356(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2291), .Q(n60[5]));
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2292), .Q(n60[6]));
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2289), .Q(n60[7]));
    or g359(n2295 ,n1436 ,n2286);
    or g360(n2294 ,n1433 ,n2287);
    or g361(n2293 ,n1430 ,n2285);
    or g362(n2292 ,n1434 ,n2282);
    or g363(n2291 ,n1435 ,n2283);
    or g364(n2290 ,n1432 ,n2288);
    or g365(n2289 ,n1431 ,n2281);
    or g366(n2288 ,n743 ,n2273);
    or g367(n2287 ,n739 ,n2277);
    or g368(n2286 ,n742 ,n2280);
    or g369(n2285 ,n737 ,n2275);
    or g370(n2284 ,n1488 ,n2278);
    or g371(n2283 ,n740 ,n2268);
    or g372(n2282 ,n738 ,n2271);
    or g373(n2281 ,n741 ,n2270);
    or g374(n2280 ,n1512 ,n2262);
    or g375(n2279 ,n1172 ,n2255);
    or g376(n2278 ,n1437 ,n2260);
    or g377(n2277 ,n1555 ,n2263);
    or g378(n2276 ,n1184 ,n2252);
    or g379(n2275 ,n1518 ,n2261);
    or g380(n2274 ,n1153 ,n2254);
    or g381(n2273 ,n1462 ,n2264);
    or g382(n2272 ,n1142 ,n2251);
    or g383(n2271 ,n1489 ,n2258);
    or g384(n2270 ,n1449 ,n2257);
    or g385(n2269 ,n1169 ,n2253);
    or g386(n2268 ,n1499 ,n2259);
    or g387(n2267 ,n1150 ,n2256);
    or g388(n2266 ,n1126 ,n2250);
    or g389(n2265 ,n1198 ,n2249);
    or g390(n2264 ,n1918 ,n2241);
    or g391(n2263 ,n1929 ,n2246);
    or g392(n2262 ,n1924 ,n2247);
    or g393(n2261 ,n1921 ,n2248);
    or g394(n2260 ,n1932 ,n2244);
    or g395(n2259 ,n1915 ,n2240);
    or g396(n2258 ,n1911 ,n2239);
    or g397(n2257 ,n1908 ,n2238);
    or g398(n2256 ,n1084 ,n2236);
    or g399(n2255 ,n1085 ,n2245);
    or g400(n2254 ,n1086 ,n2242);
    or g401(n2253 ,n1087 ,n2237);
    or g402(n2252 ,n1080 ,n2243);
    or g403(n2251 ,n1083 ,n2235);
    or g404(n2250 ,n1082 ,n2234);
    or g405(n2249 ,n1081 ,n2233);
    or g406(n2248 ,n1664 ,n2221);
    or g407(n2247 ,n1634 ,n2222);
    or g408(n2246 ,n1640 ,n2232);
    or g409(n2245 ,n1822 ,n2223);
    or g410(n2244 ,n1648 ,n2224);
    or g411(n2243 ,n1826 ,n2231);
    or g412(n2242 ,n1827 ,n2230);
    or g413(n2241 ,n1622 ,n2220);
    or g414(n2240 ,n1616 ,n2219);
    or g415(n2239 ,n1612 ,n2218);
    or g416(n2238 ,n1607 ,n2217);
    or g417(n2237 ,n1833 ,n2229);
    or g418(n2236 ,n1836 ,n2228);
    or g419(n2235 ,n1839 ,n2226);
    or g420(n2234 ,n1840 ,n2227);
    or g421(n2233 ,n1843 ,n2225);
    or g422(n2232 ,n1530 ,n2203);
    or g423(n2231 ,n1389 ,n2191);
    or g424(n2230 ,n1344 ,n2189);
    or g425(n2229 ,n1364 ,n2182);
    or g426(n2228 ,n1325 ,n2178);
    or g427(n2227 ,n1277 ,n2173);
    or g428(n2226 ,n1259 ,n2172);
    or g429(n2225 ,n1235 ,n2170);
    or g430(n2224 ,n1538 ,n2204);
    or g431(n2223 ,n1394 ,n2194);
    or g432(n2222 ,n1524 ,n2202);
    or g433(n2221 ,n1513 ,n2201);
    or g434(n2220 ,n1503 ,n2200);
    or g435(n2219 ,n1541 ,n2199);
    or g436(n2218 ,n1546 ,n2198);
    or g437(n2217 ,n1508 ,n2197);
    or g438(n2216 ,n1813 ,n2207);
    or g439(n2215 ,n1818 ,n2206);
    or g440(n2214 ,n1819 ,n2205);
    or g441(n2213 ,n1854 ,n2001);
    or g442(n2212 ,n1763 ,n2002);
    or g443(n2211 ,n1758 ,n2003);
    or g444(n2210 ,n1759 ,n2004);
    or g445(n2209 ,n1760 ,n2005);
    or g446(n2208 ,n1761 ,n2006);
    nor g447(n2207 ,n322 ,n1979);
    nor g448(n2206 ,n326 ,n1979);
    nor g449(n2205 ,n297 ,n1979);
    or g450(n2204 ,n1931 ,n1930);
    or g451(n2203 ,n1926 ,n1978);
    or g452(n2202 ,n1923 ,n1922);
    or g453(n2201 ,n1920 ,n1919);
    or g454(n2200 ,n1917 ,n1916);
    or g455(n2199 ,n1913 ,n1912);
    or g456(n2198 ,n1906 ,n1909);
    or g457(n2197 ,n1927 ,n1907);
    or g458(n2196 ,n2032 ,n1899);
    or g459(n2195 ,n2024 ,n1898);
    or g460(n2194 ,n1185 ,n1928);
    or g461(n2193 ,n2016 ,n1897);
    or g462(n2192 ,n2061 ,n1896);
    or g463(n2191 ,n1187 ,n1914);
    or g464(n2190 ,n1940 ,n1895);
    or g465(n2189 ,n1160 ,n1910);
    or g466(n2188 ,n1817 ,n1877);
    or g467(n2187 ,n1815 ,n1876);
    or g468(n2186 ,n1816 ,n1875);
    or g469(n2185 ,n1820 ,n1874);
    or g470(n2184 ,n2000 ,n1893);
    or g471(n2183 ,n1992 ,n1892);
    or g472(n2182 ,n1161 ,n1905);
    or g473(n2181 ,n1984 ,n1891);
    or g474(n2180 ,n2040 ,n1890);
    or g475(n2179 ,n2048 ,n1889);
    or g476(n2178 ,n1141 ,n1904);
    or g477(n2177 ,n2056 ,n1888);
    or g478(n2176 ,n1975 ,n1887);
    or g479(n2175 ,n1967 ,n1886);
    or g480(n2174 ,n1959 ,n1885);
    or g481(n2173 ,n1114 ,n1903);
    or g482(n2172 ,n1094 ,n1902);
    or g483(n2171 ,n1951 ,n1884);
    or g484(n2170 ,n1090 ,n1901);
    or g485(n2169 ,n1943 ,n1883);
    nor g486(n2168 ,n142 ,n1900);
    or g487(n2167 ,n1784 ,n2037);
    or g488(n2166 ,n1783 ,n2036);
    or g489(n2165 ,n1782 ,n2035);
    or g490(n2164 ,n1781 ,n2034);
    or g491(n2163 ,n1846 ,n2033);
    or g492(n2162 ,n1780 ,n2031);
    or g493(n2161 ,n1779 ,n2030);
    or g494(n2160 ,n1778 ,n2029);
    or g495(n2159 ,n1777 ,n2028);
    or g496(n2158 ,n1776 ,n2027);
    or g497(n2157 ,n1775 ,n2026);
    or g498(n2156 ,n1848 ,n2025);
    or g499(n2155 ,n1774 ,n2023);
    or g500(n2154 ,n1773 ,n2022);
    or g501(n2153 ,n1772 ,n2021);
    or g502(n2152 ,n1771 ,n2020);
    or g503(n2151 ,n1770 ,n2019);
    or g504(n2150 ,n1769 ,n2018);
    or g505(n2149 ,n1850 ,n2017);
    or g506(n2148 ,n1768 ,n2015);
    or g507(n2147 ,n1767 ,n2014);
    or g508(n2146 ,n1766 ,n2013);
    or g509(n2145 ,n1700 ,n2012);
    or g510(n2144 ,n1764 ,n2010);
    or g511(n2143 ,n1765 ,n2011);
    or g512(n2142 ,n1852 ,n2009);
    or g513(n2141 ,n1762 ,n2007);
    or g514(n2140 ,n1689 ,n1941);
    or g515(n2139 ,n1756 ,n1938);
    or g516(n2138 ,n1755 ,n1937);
    or g517(n2137 ,n1754 ,n1936);
    or g518(n2136 ,n1753 ,n1935);
    or g519(n2135 ,n1752 ,n1934);
    or g520(n2134 ,n1856 ,n1933);
    or g521(n2133 ,n1751 ,n1999);
    or g522(n2132 ,n1750 ,n1998);
    or g523(n2131 ,n1749 ,n1997);
    or g524(n2130 ,n1748 ,n1996);
    or g525(n2129 ,n1747 ,n1995);
    or g526(n2128 ,n1746 ,n1994);
    or g527(n2127 ,n1858 ,n1993);
    or g528(n2126 ,n1745 ,n1991);
    or g529(n2125 ,n1744 ,n1990);
    or g530(n2124 ,n1743 ,n1989);
    or g531(n2123 ,n1742 ,n1988);
    or g532(n2122 ,n1741 ,n1987);
    or g533(n2121 ,n1740 ,n1986);
    or g534(n2120 ,n1860 ,n1985);
    or g535(n2119 ,n1739 ,n1983);
    or g536(n2118 ,n1738 ,n1982);
    or g537(n2117 ,n1737 ,n1981);
    or g538(n2116 ,n1736 ,n1980);
    or g539(n2115 ,n1735 ,n2008);
    or g540(n2114 ,n1734 ,n2038);
    or g541(n2113 ,n1862 ,n2039);
    or g542(n2112 ,n1733 ,n2041);
    or g543(n2111 ,n1732 ,n2042);
    or g544(n2110 ,n1731 ,n2043);
    or g545(n2109 ,n1730 ,n2044);
    or g546(n2108 ,n1729 ,n2045);
    or g547(n2107 ,n1728 ,n2046);
    or g548(n2106 ,n1864 ,n2047);
    or g549(n2105 ,n1727 ,n2049);
    or g550(n2104 ,n1726 ,n2050);
    or g551(n2103 ,n1725 ,n2051);
    or g552(n2102 ,n1724 ,n2052);
    or g553(n2101 ,n1723 ,n2053);
    or g554(n2100 ,n1722 ,n2054);
    or g555(n2099 ,n1866 ,n2055);
    or g556(n2098 ,n1721 ,n2057);
    or g557(n2097 ,n1720 ,n2058);
    or g558(n2096 ,n1719 ,n2059);
    or g559(n2095 ,n1718 ,n2060);
    or g560(n2094 ,n1717 ,n1925);
    or g561(n2093 ,n1716 ,n1977);
    or g562(n2092 ,n1868 ,n1976);
    or g563(n2091 ,n1715 ,n1974);
    or g564(n2090 ,n1714 ,n1973);
    or g565(n2089 ,n1713 ,n1972);
    or g566(n2088 ,n1712 ,n1971);
    or g567(n2087 ,n1711 ,n1970);
    or g568(n2086 ,n1710 ,n1968);
    or g569(n2085 ,n1870 ,n1969);
    or g570(n2084 ,n1709 ,n1966);
    or g571(n2083 ,n1708 ,n1965);
    or g572(n2082 ,n1707 ,n1964);
    or g573(n2081 ,n1706 ,n1963);
    or g574(n2080 ,n1705 ,n1962);
    or g575(n2079 ,n1704 ,n1961);
    or g576(n2078 ,n1872 ,n1960);
    or g577(n2077 ,n1703 ,n1958);
    or g578(n2076 ,n1702 ,n1957);
    or g579(n2075 ,n1701 ,n1956);
    or g580(n2074 ,n1699 ,n1955);
    or g581(n2073 ,n1698 ,n1954);
    or g582(n2072 ,n1697 ,n1953);
    or g583(n2071 ,n1788 ,n1952);
    or g584(n2070 ,n1696 ,n1950);
    or g585(n2069 ,n1695 ,n1949);
    or g586(n2068 ,n1694 ,n1948);
    or g587(n2067 ,n1693 ,n1947);
    or g588(n2066 ,n1692 ,n1946);
    or g589(n2065 ,n1691 ,n1945);
    or g590(n2064 ,n1786 ,n1944);
    or g591(n2063 ,n1690 ,n1942);
    or g592(n2062 ,n1757 ,n1939);
    nor g593(n2061 ,n379 ,n1792);
    nor g594(n2060 ,n418 ,n1799);
    nor g595(n2059 ,n485 ,n1799);
    nor g596(n2058 ,n398 ,n1799);
    nor g597(n2057 ,n424 ,n1799);
    nor g598(n2056 ,n251 ,n1799);
    nor g599(n2055 ,n260 ,n1798);
    nor g600(n2054 ,n461 ,n1798);
    nor g601(n2053 ,n202 ,n1798);
    nor g602(n2052 ,n430 ,n1798);
    nor g603(n2051 ,n405 ,n1798);
    nor g604(n2050 ,n425 ,n1798);
    nor g605(n2049 ,n438 ,n1798);
    nor g606(n2048 ,n195 ,n1798);
    nor g607(n2047 ,n183 ,n1797);
    nor g608(n2046 ,n370 ,n1797);
    nor g609(n2045 ,n275 ,n1797);
    nor g610(n2044 ,n292 ,n1797);
    nor g611(n2043 ,n472 ,n1797);
    nor g612(n2042 ,n287 ,n1797);
    nor g613(n2041 ,n381 ,n1797);
    nor g614(n2040 ,n356 ,n1797);
    nor g615(n2039 ,n230 ,n1796);
    nor g616(n2038 ,n384 ,n1796);
    nor g617(n2037 ,n281 ,n1793);
    nor g618(n2036 ,n276 ,n1793);
    nor g619(n2035 ,n469 ,n1793);
    nor g620(n2034 ,n368 ,n1793);
    nor g621(n2033 ,n177 ,n1793);
    nor g622(n2032 ,n432 ,n1804);
    nor g623(n2031 ,n477 ,n1804);
    nor g624(n2030 ,n282 ,n1804);
    nor g625(n2029 ,n182 ,n1804);
    nor g626(n2028 ,n491 ,n1804);
    nor g627(n2027 ,n209 ,n1804);
    nor g628(n2026 ,n436 ,n1804);
    nor g629(n2025 ,n402 ,n1804);
    nor g630(n2024 ,n273 ,n1790);
    nor g631(n2023 ,n396 ,n1790);
    nor g632(n2022 ,n219 ,n1790);
    nor g633(n2021 ,n363 ,n1790);
    nor g634(n2020 ,n193 ,n1790);
    nor g635(n2019 ,n502 ,n1790);
    nor g636(n2018 ,n270 ,n1790);
    nor g637(n2017 ,n374 ,n1790);
    nor g638(n2016 ,n476 ,n1791);
    nor g639(n2015 ,n176 ,n1791);
    nor g640(n2014 ,n495 ,n1791);
    nor g641(n2013 ,n474 ,n1791);
    nor g642(n2012 ,n191 ,n1791);
    nor g643(n2011 ,n203 ,n1791);
    nor g644(n2010 ,n284 ,n1791);
    nor g645(n2009 ,n205 ,n1791);
    nor g646(n2008 ,n408 ,n1796);
    nor g647(n2007 ,n214 ,n1792);
    nor g648(n2006 ,n247 ,n1792);
    nor g649(n2005 ,n475 ,n1792);
    nor g650(n2004 ,n391 ,n1792);
    nor g651(n2003 ,n395 ,n1792);
    nor g652(n2002 ,n295 ,n1792);
    nor g653(n2001 ,n488 ,n1792);
    nor g654(n2000 ,n185 ,n1794);
    nor g655(n1999 ,n479 ,n1794);
    nor g656(n1998 ,n208 ,n1794);
    nor g657(n1997 ,n468 ,n1794);
    nor g658(n1996 ,n421 ,n1794);
    nor g659(n1995 ,n239 ,n1794);
    nor g660(n1994 ,n234 ,n1794);
    nor g661(n1993 ,n416 ,n1794);
    nor g662(n1992 ,n400 ,n1795);
    nor g663(n1991 ,n393 ,n1795);
    nor g664(n1990 ,n357 ,n1795);
    nor g665(n1989 ,n390 ,n1795);
    nor g666(n1988 ,n245 ,n1795);
    nor g667(n1987 ,n389 ,n1795);
    nor g668(n1986 ,n434 ,n1795);
    nor g669(n1985 ,n236 ,n1795);
    nor g670(n1984 ,n437 ,n1796);
    nor g671(n1983 ,n371 ,n1796);
    nor g672(n1982 ,n417 ,n1796);
    nor g673(n1981 ,n361 ,n1796);
    nor g674(n1980 ,n453 ,n1796);
    or g675(n1978 ,n1637 ,n1636);
    nor g676(n1977 ,n222 ,n1799);
    nor g677(n1976 ,n442 ,n1799);
    nor g678(n1975 ,n497 ,n1800);
    nor g679(n1974 ,n428 ,n1800);
    nor g680(n1973 ,n467 ,n1800);
    nor g681(n1972 ,n509 ,n1800);
    nor g682(n1971 ,n455 ,n1800);
    nor g683(n1970 ,n466 ,n1800);
    nor g684(n1969 ,n204 ,n1800);
    nor g685(n1968 ,n358 ,n1800);
    nor g686(n1967 ,n464 ,n1801);
    nor g687(n1966 ,n226 ,n1801);
    nor g688(n1965 ,n447 ,n1801);
    nor g689(n1964 ,n382 ,n1801);
    nor g690(n1963 ,n470 ,n1801);
    nor g691(n1962 ,n478 ,n1801);
    nor g692(n1961 ,n244 ,n1801);
    nor g693(n1960 ,n354 ,n1801);
    nor g694(n1959 ,n175 ,n1802);
    nor g695(n1958 ,n268 ,n1802);
    nor g696(n1957 ,n257 ,n1802);
    nor g697(n1956 ,n217 ,n1802);
    nor g698(n1955 ,n378 ,n1802);
    nor g699(n1954 ,n406 ,n1802);
    nor g700(n1953 ,n232 ,n1802);
    nor g701(n1952 ,n254 ,n1802);
    nor g702(n1951 ,n197 ,n1803);
    nor g703(n1950 ,n221 ,n1803);
    nor g704(n1949 ,n501 ,n1803);
    nor g705(n1948 ,n459 ,n1803);
    nor g706(n1947 ,n243 ,n1803);
    nor g707(n1946 ,n465 ,n1803);
    nor g708(n1945 ,n510 ,n1803);
    nor g709(n1944 ,n365 ,n1803);
    nor g710(n1943 ,n503 ,n1793);
    nor g711(n1942 ,n194 ,n1793);
    nor g712(n1941 ,n484 ,n1793);
    nor g713(n1940 ,n355 ,n1789);
    nor g714(n1939 ,n399 ,n1789);
    nor g715(n1938 ,n376 ,n1789);
    nor g716(n1937 ,n218 ,n1789);
    nor g717(n1936 ,n407 ,n1789);
    nor g718(n1935 ,n367 ,n1789);
    nor g719(n1934 ,n494 ,n1789);
    nor g720(n1933 ,n360 ,n1789);
    or g721(n1932 ,n1650 ,n1649);
    or g722(n1931 ,n1647 ,n1646);
    or g723(n1930 ,n1645 ,n1644);
    or g724(n1929 ,n1641 ,n1657);
    or g725(n1928 ,n1824 ,n1825);
    or g726(n1927 ,n1606 ,n1655);
    or g727(n1926 ,n1639 ,n1638);
    nor g728(n1925 ,n493 ,n1799);
    or g729(n1924 ,n1666 ,n1635);
    or g730(n1923 ,n1633 ,n1632);
    or g731(n1922 ,n1669 ,n1631);
    or g732(n1921 ,n1667 ,n1629);
    or g733(n1920 ,n1665 ,n1627);
    or g734(n1919 ,n1626 ,n1625);
    or g735(n1918 ,n1624 ,n1623);
    or g736(n1917 ,n1621 ,n1620);
    or g737(n1916 ,n1611 ,n1619);
    or g738(n1915 ,n1618 ,n1617);
    or g739(n1914 ,n1831 ,n1830);
    or g740(n1913 ,n1654 ,n1615);
    or g741(n1912 ,n1668 ,n1614);
    or g742(n1911 ,n1643 ,n1613);
    or g743(n1910 ,n1828 ,n1829);
    or g744(n1909 ,n1662 ,n1628);
    or g745(n1908 ,n1609 ,n1608);
    or g746(n1907 ,n1630 ,n1656);
    or g747(n1906 ,n1610 ,n1642);
    or g748(n1905 ,n1834 ,n1835);
    or g749(n1904 ,n1837 ,n1838);
    or g750(n1903 ,n1841 ,n1842);
    or g751(n1902 ,n1844 ,n1823);
    or g752(n1901 ,n1845 ,n1821);
    nor g753(n1900 ,n1812 ,n1686);
    or g754(n1899 ,n147 ,n1847);
    or g755(n1898 ,n146 ,n1849);
    or g756(n1897 ,n145 ,n1851);
    or g757(n1896 ,n147 ,n1853);
    or g758(n1895 ,n146 ,n1855);
    nor g759(n1894 ,n143 ,n1670);
    or g760(n1893 ,n145 ,n1857);
    or g761(n1892 ,n146 ,n1859);
    or g762(n1891 ,n147 ,n1861);
    or g763(n1890 ,n141 ,n1863);
    or g764(n1889 ,n141 ,n1865);
    or g765(n1888 ,n144 ,n1867);
    or g766(n1887 ,n141 ,n1869);
    or g767(n1886 ,n147 ,n1871);
    or g768(n1885 ,n146 ,n1873);
    or g769(n1884 ,n144 ,n1787);
    or g770(n1883 ,n144 ,n1785);
    or g771(n1882 ,n728 ,n1805);
    or g772(n1881 ,n744 ,n1806);
    or g773(n1880 ,n727 ,n1807);
    or g774(n1879 ,n546 ,n1832);
    or g775(n1878 ,n1814 ,n1687);
    or g776(n1877 ,n610 ,n1808);
    or g777(n1876 ,n607 ,n1809);
    or g778(n1875 ,n609 ,n1810);
    or g779(n1874 ,n608 ,n1811);
    or g780(n1979 ,n995 ,n1789);
    nor g781(n1873 ,n2296 ,n1588);
    nor g782(n1872 ,n151 ,n1572);
    nor g783(n1871 ,n2296 ,n1572);
    nor g784(n1870 ,n151 ,n1584);
    nor g785(n1869 ,n2296 ,n1584);
    nor g786(n1868 ,n151 ,n1582);
    nor g787(n1867 ,n2296 ,n1582);
    nor g788(n1866 ,n151 ,n1580);
    nor g789(n1865 ,n2296 ,n1580);
    nor g790(n1864 ,n151 ,n1578);
    nor g791(n1863 ,n2296 ,n1578);
    nor g792(n1862 ,n151 ,n1598);
    nor g793(n1861 ,n2296 ,n1598);
    nor g794(n1860 ,n151 ,n1576);
    nor g795(n1859 ,n2296 ,n1576);
    nor g796(n1858 ,n151 ,n1594);
    nor g797(n1857 ,n2296 ,n1594);
    nor g798(n1856 ,n151 ,n1590);
    nor g799(n1855 ,n2296 ,n1590);
    nor g800(n1854 ,n151 ,n1600);
    nor g801(n1853 ,n2296 ,n1600);
    nor g802(n1852 ,n151 ,n1592);
    nor g803(n1851 ,n2296 ,n1592);
    nor g804(n1850 ,n151 ,n1586);
    nor g805(n1849 ,n2296 ,n1586);
    nor g806(n1848 ,n151 ,n1602);
    nor g807(n1847 ,n2296 ,n1602);
    nor g808(n1846 ,n151 ,n1574);
    or g809(n1845 ,n1231 ,n1228);
    or g810(n1844 ,n1236 ,n1233);
    or g811(n1843 ,n1243 ,n1241);
    or g812(n1842 ,n1260 ,n1256);
    or g813(n1841 ,n1268 ,n1265);
    or g814(n1840 ,n1287 ,n1285);
    or g815(n1839 ,n1294 ,n1289);
    or g816(n1838 ,n1303 ,n1299);
    or g817(n1837 ,n1313 ,n1308);
    or g818(n1836 ,n1330 ,n1329);
    or g819(n1835 ,n1347 ,n1342);
    or g820(n1834 ,n1356 ,n1348);
    or g821(n1833 ,n1370 ,n1369);
    nor g822(n1832 ,n726 ,n1603);
    or g823(n1831 ,n1391 ,n1384);
    or g824(n1830 ,n1380 ,n1376);
    or g825(n1829 ,n1385 ,n1382);
    or g826(n1828 ,n1392 ,n1386);
    or g827(n1827 ,n1383 ,n1388);
    or g828(n1826 ,n1254 ,n1320);
    or g829(n1825 ,n1258 ,n1279);
    or g830(n1824 ,n1393 ,n1250);
    or g831(n1823 ,n1292 ,n1358);
    or g832(n1822 ,n1367 ,n1395);
    or g833(n1821 ,n1403 ,n1399);
    nor g834(n1820 ,n163 ,n1411);
    nor g835(n1819 ,n166 ,n1603);
    nor g836(n1818 ,n334 ,n1603);
    nor g837(n1817 ,n169 ,n1411);
    nor g838(n1816 ,n345 ,n1411);
    nor g839(n1815 ,n171 ,n1411);
    nor g840(n1814 ,n347 ,n1411);
    nor g841(n1813 ,n342 ,n1603);
    nor g842(n1812 ,n403 ,n1413);
    nor g843(n1811 ,n301 ,n1604);
    nor g844(n1810 ,n307 ,n1604);
    nor g845(n1809 ,n309 ,n1604);
    nor g846(n1808 ,n311 ,n1604);
    nor g847(n1807 ,n302 ,n1605);
    nor g848(n1806 ,n314 ,n1605);
    nor g849(n1805 ,n313 ,n1605);
    nor g850(n1788 ,n151 ,n1588);
    nor g851(n1787 ,n2296 ,n1596);
    nor g852(n1786 ,n151 ,n1596);
    nor g853(n1785 ,n2296 ,n1574);
    nor g854(n1784 ,n328 ,n1574);
    nor g855(n1783 ,n327 ,n1574);
    nor g856(n1782 ,n329 ,n1574);
    nor g857(n1781 ,n150 ,n1574);
    nor g858(n1780 ,n149 ,n1602);
    nor g859(n1779 ,n148 ,n1602);
    nor g860(n1778 ,n328 ,n1602);
    nor g861(n1777 ,n327 ,n1602);
    nor g862(n1776 ,n329 ,n1602);
    nor g863(n1775 ,n150 ,n1602);
    nor g864(n1774 ,n149 ,n1586);
    nor g865(n1773 ,n148 ,n1586);
    nor g866(n1772 ,n328 ,n1586);
    nor g867(n1771 ,n327 ,n1586);
    nor g868(n1770 ,n329 ,n1586);
    nor g869(n1769 ,n150 ,n1586);
    nor g870(n1768 ,n149 ,n1592);
    nor g871(n1767 ,n148 ,n1592);
    nor g872(n1766 ,n328 ,n1592);
    nor g873(n1765 ,n329 ,n1592);
    nor g874(n1764 ,n150 ,n1592);
    nor g875(n1763 ,n150 ,n1600);
    nor g876(n1762 ,n149 ,n1600);
    nor g877(n1761 ,n148 ,n1600);
    nor g878(n1760 ,n328 ,n1600);
    nor g879(n1759 ,n327 ,n1600);
    nor g880(n1758 ,n329 ,n1600);
    nor g881(n1757 ,n149 ,n1590);
    nor g882(n1756 ,n148 ,n1590);
    nor g883(n1755 ,n328 ,n1590);
    nor g884(n1754 ,n327 ,n1590);
    nor g885(n1753 ,n329 ,n1590);
    nor g886(n1752 ,n150 ,n1590);
    nor g887(n1751 ,n149 ,n1594);
    nor g888(n1750 ,n148 ,n1594);
    nor g889(n1749 ,n328 ,n1594);
    nor g890(n1748 ,n327 ,n1594);
    nor g891(n1747 ,n329 ,n1594);
    nor g892(n1746 ,n150 ,n1594);
    nor g893(n1745 ,n149 ,n1576);
    nor g894(n1744 ,n148 ,n1576);
    nor g895(n1743 ,n328 ,n1576);
    nor g896(n1742 ,n327 ,n1576);
    nor g897(n1741 ,n329 ,n1576);
    nor g898(n1740 ,n150 ,n1576);
    nor g899(n1739 ,n149 ,n1598);
    nor g900(n1738 ,n148 ,n1598);
    nor g901(n1737 ,n328 ,n1598);
    nor g902(n1736 ,n327 ,n1598);
    nor g903(n1735 ,n329 ,n1598);
    nor g904(n1734 ,n150 ,n1598);
    nor g905(n1733 ,n149 ,n1578);
    nor g906(n1732 ,n148 ,n1578);
    nor g907(n1731 ,n328 ,n1578);
    nor g908(n1730 ,n327 ,n1578);
    nor g909(n1729 ,n329 ,n1578);
    nor g910(n1728 ,n150 ,n1578);
    nor g911(n1727 ,n149 ,n1580);
    nor g912(n1726 ,n148 ,n1580);
    nor g913(n1725 ,n328 ,n1580);
    nor g914(n1724 ,n327 ,n1580);
    nor g915(n1723 ,n329 ,n1580);
    nor g916(n1722 ,n150 ,n1580);
    nor g917(n1721 ,n149 ,n1582);
    nor g918(n1720 ,n148 ,n1582);
    nor g919(n1719 ,n328 ,n1582);
    nor g920(n1718 ,n327 ,n1582);
    nor g921(n1717 ,n329 ,n1582);
    nor g922(n1716 ,n150 ,n1582);
    nor g923(n1715 ,n149 ,n1584);
    nor g924(n1714 ,n148 ,n1584);
    nor g925(n1713 ,n328 ,n1584);
    nor g926(n1712 ,n327 ,n1584);
    nor g927(n1711 ,n329 ,n1584);
    nor g928(n1710 ,n150 ,n1584);
    nor g929(n1709 ,n149 ,n1572);
    nor g930(n1708 ,n148 ,n1572);
    nor g931(n1707 ,n328 ,n1572);
    nor g932(n1706 ,n327 ,n1572);
    nor g933(n1705 ,n329 ,n1572);
    nor g934(n1704 ,n150 ,n1572);
    nor g935(n1703 ,n149 ,n1588);
    nor g936(n1702 ,n148 ,n1588);
    nor g937(n1701 ,n328 ,n1588);
    nor g938(n1700 ,n327 ,n1592);
    nor g939(n1699 ,n327 ,n1588);
    nor g940(n1698 ,n329 ,n1588);
    nor g941(n1697 ,n150 ,n1588);
    nor g942(n1696 ,n149 ,n1596);
    nor g943(n1695 ,n148 ,n1596);
    nor g944(n1694 ,n328 ,n1596);
    nor g945(n1693 ,n327 ,n1596);
    nor g946(n1692 ,n329 ,n1596);
    nor g947(n1691 ,n150 ,n1596);
    nor g948(n1690 ,n149 ,n1574);
    nor g949(n1689 ,n148 ,n1574);
    or g950(n1688 ,n928 ,n1408);
    nor g951(n1687 ,n529 ,n1410);
    nor g952(n1686 ,n528 ,n1412);
    or g953(n1685 ,n859 ,n1419);
    or g954(n1684 ,n851 ,n1420);
    or g955(n1683 ,n845 ,n1421);
    or g956(n1682 ,n1036 ,n1423);
    or g957(n1681 ,n834 ,n1424);
    or g958(n1680 ,n1019 ,n1425);
    or g959(n1679 ,n1011 ,n1426);
    or g960(n1678 ,n868 ,n1427);
    or g961(n1677 ,n866 ,n1479);
    or g962(n1676 ,n961 ,n1564);
    or g963(n1675 ,n955 ,n1565);
    or g964(n1674 ,n798 ,n1566);
    or g965(n1673 ,n876 ,n1567);
    or g966(n1672 ,n1072 ,n1568);
    or g967(n1671 ,n1032 ,n1569);
    xor g968(n1670 ,n995 ,n38[0]);
    or g969(n1669 ,n1520 ,n1521);
    or g970(n1668 ,n1454 ,n1491);
    or g971(n1667 ,n1450 ,n1517);
    or g972(n1666 ,n1526 ,n1444);
    or g973(n1665 ,n1452 ,n1456);
    or g974(n1664 ,n1453 ,n1514);
    or g975(n1663 ,n1428 ,n1422);
    or g976(n1662 ,n1483 ,n1457);
    or g977(n1661 ,n1429 ,n1416);
    or g978(n1660 ,n623 ,n1558);
    or g979(n1659 ,n622 ,n1559);
    or g980(n1658 ,n618 ,n1560);
    or g981(n1657 ,n1531 ,n1202);
    or g982(n1656 ,n1472 ,n1441);
    or g983(n1655 ,n1475 ,n1570);
    or g984(n1654 ,n1493 ,n1465);
    or g985(n1653 ,n1221 ,n1563);
    or g986(n1652 ,n923 ,n1562);
    or g987(n1651 ,n1224 ,n1561);
    or g988(n1650 ,n1502 ,n1543);
    or g989(n1649 ,n1542 ,n1208);
    or g990(n1648 ,n1540 ,n1539);
    or g991(n1647 ,n1552 ,n1537);
    or g992(n1646 ,n1536 ,n1535);
    or g993(n1645 ,n1451 ,n1534);
    or g994(n1644 ,n1533 ,n1532);
    or g995(n1643 ,n1468 ,n1553);
    or g996(n1642 ,n1484 ,n1445);
    or g997(n1641 ,n1554 ,n1485);
    or g998(n1640 ,n1464 ,n1515);
    or g999(n1639 ,n1529 ,n1557);
    or g1000(n1638 ,n1547 ,n1527);
    or g1001(n1637 ,n1470 ,n1492);
    or g1002(n1636 ,n1548 ,n1528);
    or g1003(n1635 ,n1438 ,n1210);
    or g1004(n1634 ,n1525 ,n1439);
    or g1005(n1633 ,n1442 ,n1447);
    or g1006(n1632 ,n1522 ,n1446);
    or g1007(n1631 ,n1448 ,n1519);
    or g1008(n1630 ,n1473 ,n1474);
    or g1009(n1629 ,n1516 ,n1125);
    or g1010(n1628 ,n1509 ,n1481);
    or g1011(n1627 ,n1511 ,n1550);
    or g1012(n1626 ,n1461 ,n1458);
    or g1013(n1625 ,n1510 ,n1459);
    or g1014(n1624 ,n1506 ,n1463);
    or g1015(n1623 ,n1505 ,n1193);
    or g1016(n1622 ,n1504 ,n1495);
    or g1017(n1621 ,n1471 ,n1494);
    or g1018(n1620 ,n1486 ,n1482);
    or g1019(n1619 ,n1500 ,n1498);
    or g1020(n1618 ,n1440 ,n1523);
    or g1021(n1617 ,n1497 ,n1186);
    or g1022(n1616 ,n1496 ,n1544);
    or g1023(n1615 ,n1551 ,n1455);
    or g1024(n1614 ,n1490 ,n1556);
    or g1025(n1613 ,n1443 ,n1122);
    or g1026(n1612 ,n1477 ,n1469);
    or g1027(n1611 ,n1501 ,n1487);
    or g1028(n1610 ,n1460 ,n1549);
    or g1029(n1609 ,n1466 ,n1480);
    or g1030(n1608 ,n1545 ,n1199);
    or g1031(n1607 ,n1478 ,n1467);
    or g1032(n1606 ,n1476 ,n1507);
    or g1033(n1804 ,n147 ,n1601);
    or g1034(n1803 ,n147 ,n1595);
    or g1035(n1802 ,n145 ,n1587);
    or g1036(n1801 ,n141 ,n1571);
    or g1037(n1800 ,n141 ,n1583);
    or g1038(n1799 ,n141 ,n1581);
    or g1039(n1798 ,n147 ,n1579);
    or g1040(n1797 ,n146 ,n1577);
    or g1041(n1796 ,n145 ,n1597);
    or g1042(n1795 ,n146 ,n1575);
    or g1043(n1794 ,n146 ,n1593);
    or g1044(n1793 ,n146 ,n1573);
    or g1045(n1792 ,n145 ,n1599);
    or g1046(n1791 ,n145 ,n1591);
    or g1047(n1790 ,n145 ,n1585);
    or g1048(n1789 ,n147 ,n1589);
    not g1049(n1602 ,n1601);
    not g1050(n1600 ,n1599);
    not g1051(n1598 ,n1597);
    not g1052(n1596 ,n1595);
    not g1053(n1594 ,n1593);
    not g1054(n1592 ,n1591);
    not g1055(n1590 ,n1589);
    not g1056(n1588 ,n1587);
    not g1057(n1586 ,n1585);
    not g1058(n1584 ,n1583);
    not g1059(n1582 ,n1581);
    not g1060(n1580 ,n1579);
    not g1061(n1578 ,n1577);
    not g1062(n1576 ,n1575);
    not g1063(n1574 ,n1573);
    not g1064(n1572 ,n1571);
    nor g1065(n1570 ,n255 ,n993);
    or g1066(n1569 ,n147 ,n839);
    or g1067(n1568 ,n147 ,n797);
    or g1068(n1567 ,n147 ,n1070);
    or g1069(n1566 ,n145 ,n1062);
    or g1070(n1565 ,n145 ,n878);
    or g1071(n1564 ,n145 ,n807);
    nor g1072(n1563 ,n321 ,n1001);
    nor g1073(n1562 ,n310 ,n1001);
    nor g1074(n1561 ,n304 ,n1001);
    nor g1075(n1560 ,n320 ,n1004);
    nor g1076(n1559 ,n308 ,n1004);
    nor g1077(n1558 ,n325 ,n1004);
    nor g1078(n1557 ,n199 ,n980);
    nor g1079(n1556 ,n263 ,n990);
    nor g1080(n1555 ,n454 ,n984);
    nor g1081(n1554 ,n364 ,n985);
    nor g1082(n1553 ,n252 ,n994);
    nor g1083(n1552 ,n266 ,n982);
    nor g1084(n1551 ,n452 ,n988);
    nor g1085(n1550 ,n267 ,n993);
    nor g1086(n1549 ,n264 ,n980);
    nor g1087(n1548 ,n498 ,n983);
    nor g1088(n1547 ,n274 ,n988);
    nor g1089(n1546 ,n269 ,n989);
    nor g1090(n1545 ,n413 ,n992);
    nor g1091(n1544 ,n486 ,n986);
    nor g1092(n1543 ,n483 ,n994);
    nor g1093(n1542 ,n256 ,n992);
    nor g1094(n1541 ,n496 ,n989);
    nor g1095(n1540 ,n435 ,n987);
    nor g1096(n1539 ,n415 ,n986);
    nor g1097(n1538 ,n431 ,n989);
    nor g1098(n1537 ,n482 ,n980);
    nor g1099(n1536 ,n352 ,n988);
    nor g1100(n1535 ,n288 ,n993);
    nor g1101(n1534 ,n471 ,n991);
    nor g1102(n1533 ,n190 ,n983);
    nor g1103(n1532 ,n450 ,n990);
    nor g1104(n1531 ,n505 ,n992);
    nor g1105(n1530 ,n242 ,n989);
    nor g1106(n1529 ,n186 ,n982);
    nor g1107(n1528 ,n283 ,n990);
    nor g1108(n1527 ,n427 ,n993);
    nor g1109(n1526 ,n362 ,n985);
    nor g1110(n1525 ,n184 ,n987);
    nor g1111(n1524 ,n253 ,n989);
    nor g1112(n1523 ,n248 ,n994);
    nor g1113(n1522 ,n401 ,n988);
    nor g1114(n1521 ,n448 ,n991);
    nor g1115(n1520 ,n380 ,n981);
    nor g1116(n1519 ,n353 ,n990);
    nor g1117(n1518 ,n201 ,n984);
    nor g1118(n1517 ,n473 ,n994);
    nor g1119(n1516 ,n508 ,n992);
    nor g1120(n1515 ,n359 ,n986);
    nor g1121(n1514 ,n290 ,n986);
    nor g1122(n1513 ,n444 ,n989);
    nor g1123(n1512 ,n426 ,n984);
    nor g1124(n1511 ,n237 ,n988);
    nor g1125(n1510 ,n278 ,n983);
    nor g1126(n1509 ,n422 ,n983);
    nor g1127(n1508 ,n246 ,n989);
    nor g1128(n1507 ,n259 ,n980);
    nor g1129(n1506 ,n397 ,n985);
    nor g1130(n1505 ,n507 ,n992);
    nor g1131(n1504 ,n272 ,n987);
    nor g1132(n1503 ,n225 ,n989);
    nor g1133(n1502 ,n500 ,n985);
    nor g1134(n1501 ,n439 ,n981);
    nor g1135(n1500 ,n423 ,n983);
    nor g1136(n1499 ,n443 ,n984);
    nor g1137(n1498 ,n241 ,n990);
    nor g1138(n1497 ,n265 ,n992);
    nor g1139(n1496 ,n377 ,n987);
    nor g1140(n1495 ,n210 ,n986);
    nor g1141(n1494 ,n258 ,n980);
    nor g1142(n1493 ,n412 ,n982);
    nor g1143(n1492 ,n277 ,n991);
    nor g1144(n1491 ,n433 ,n991);
    nor g1145(n1490 ,n215 ,n983);
    nor g1146(n1489 ,n386 ,n984);
    nor g1147(n1488 ,n212 ,n984);
    nor g1148(n1487 ,n206 ,n991);
    nor g1149(n1486 ,n233 ,n988);
    nor g1150(n1485 ,n286 ,n994);
    nor g1151(n1484 ,n404 ,n988);
    nor g1152(n1483 ,n228 ,n981);
    nor g1153(n1482 ,n285 ,n993);
    nor g1154(n1481 ,n366 ,n990);
    nor g1155(n1480 ,n449 ,n994);
    or g1156(n1479 ,n147 ,n1074);
    nor g1157(n1478 ,n411 ,n987);
    nor g1158(n1477 ,n445 ,n987);
    nor g1159(n1476 ,n289 ,n982);
    nor g1160(n1475 ,n410 ,n988);
    nor g1161(n1474 ,n446 ,n991);
    nor g1162(n1473 ,n373 ,n981);
    nor g1163(n1472 ,n487 ,n983);
    nor g1164(n1471 ,n492 ,n982);
    nor g1165(n1470 ,n262 ,n981);
    nor g1166(n1469 ,n207 ,n986);
    nor g1167(n1468 ,n383 ,n985);
    nor g1168(n1467 ,n174 ,n986);
    nor g1169(n1466 ,n504 ,n985);
    nor g1170(n1465 ,n490 ,n980);
    nor g1171(n1464 ,n220 ,n987);
    nor g1172(n1463 ,n414 ,n994);
    nor g1173(n1462 ,n240 ,n984);
    nor g1174(n1461 ,n489 ,n981);
    nor g1175(n1460 ,n261 ,n982);
    nor g1176(n1459 ,n481 ,n990);
    nor g1177(n1458 ,n294 ,n991);
    nor g1178(n1457 ,n271 ,n991);
    nor g1179(n1456 ,n238 ,n980);
    nor g1180(n1455 ,n213 ,n993);
    nor g1181(n1454 ,n457 ,n981);
    nor g1182(n1453 ,n419 ,n987);
    nor g1183(n1452 ,n480 ,n982);
    nor g1184(n1451 ,n499 ,n981);
    nor g1185(n1450 ,n293 ,n985);
    nor g1186(n1449 ,n280 ,n984);
    nor g1187(n1448 ,n506 ,n983);
    nor g1188(n1447 ,n394 ,n980);
    nor g1189(n1446 ,n372 ,n993);
    nor g1190(n1445 ,n181 ,n993);
    nor g1191(n1444 ,n231 ,n994);
    nor g1192(n1443 ,n463 ,n992);
    nor g1193(n1442 ,n429 ,n982);
    nor g1194(n1441 ,n249 ,n990);
    nor g1195(n1440 ,n387 ,n985);
    nor g1196(n1439 ,n224 ,n986);
    nor g1197(n1438 ,n250 ,n992);
    nor g1198(n1437 ,n223 ,n979);
    nor g1199(n1436 ,n458 ,n979);
    nor g1200(n1435 ,n420 ,n979);
    nor g1201(n1434 ,n180 ,n979);
    nor g1202(n1433 ,n440 ,n979);
    nor g1203(n1432 ,n179 ,n979);
    nor g1204(n1431 ,n369 ,n979);
    nor g1205(n1430 ,n392 ,n979);
    nor g1206(n1429 ,n161 ,n1003);
    nor g1207(n1428 ,n160 ,n1003);
    or g1208(n1427 ,n146 ,n1115);
    or g1209(n1426 ,n146 ,n823);
    or g1210(n1425 ,n145 ,n828);
    or g1211(n1424 ,n145 ,n1027);
    or g1212(n1423 ,n144 ,n838);
    nor g1213(n1422 ,n643 ,n924);
    or g1214(n1421 ,n144 ,n1043);
    or g1215(n1420 ,n146 ,n1052);
    or g1216(n1419 ,n141 ,n1061);
    or g1217(n1418 ,n1218 ,n918);
    or g1218(n1417 ,n1217 ,n920);
    nor g1219(n1416 ,n597 ,n1002);
    or g1220(n1415 ,n922 ,n977);
    or g1221(n1414 ,n1219 ,n919);
    or g1222(n1605 ,n587 ,n978);
    or g1223(n1604 ,n146 ,n995);
    or g1224(n1603 ,n146 ,n996);
    nor g1225(n1601 ,n771 ,n998);
    nor g1226(n1599 ,n773 ,n997);
    nor g1227(n1597 ,n720 ,n998);
    nor g1228(n1595 ,n771 ,n999);
    nor g1229(n1593 ,n720 ,n999);
    nor g1230(n1591 ,n771 ,n1000);
    nor g1231(n1589 ,n771 ,n997);
    nor g1232(n1587 ,n773 ,n999);
    nor g1233(n1585 ,n773 ,n1000);
    nor g1234(n1583 ,n720 ,n997);
    nor g1235(n1581 ,n719 ,n1000);
    nor g1236(n1579 ,n720 ,n1000);
    nor g1237(n1577 ,n719 ,n998);
    nor g1238(n1575 ,n719 ,n999);
    nor g1239(n1573 ,n773 ,n998);
    nor g1240(n1571 ,n719 ,n997);
    not g1241(n1413 ,n1412);
    not g1242(n1411 ,n1410);
    or g1243(n1409 ,n781 ,n927);
    or g1244(n1408 ,n147 ,n776);
    or g1245(n1407 ,n777 ,n1079);
    or g1246(n1406 ,n730 ,n1223);
    or g1247(n1405 ,n778 ,n1078);
    or g1248(n1404 ,n779 ,n1077);
    or g1249(n1403 ,n1215 ,n1091);
    or g1250(n1402 ,n780 ,n1025);
    or g1251(n1401 ,n783 ,n1014);
    or g1252(n1400 ,n1216 ,n915);
    or g1253(n1399 ,n1104 ,n1214);
    or g1254(n1398 ,n731 ,n1222);
    or g1255(n1397 ,n901 ,n950);
    or g1256(n1396 ,n688 ,n926);
    or g1257(n1395 ,n1195 ,n1203);
    or g1258(n1394 ,n1099 ,n1205);
    or g1259(n1393 ,n1175 ,n1173);
    or g1260(n1392 ,n1190 ,n1201);
    or g1261(n1391 ,n1135 ,n1181);
    or g1262(n1390 ,n887 ,n1071);
    or g1263(n1389 ,n1149 ,n1144);
    or g1264(n1388 ,n1197 ,n1117);
    or g1265(n1387 ,n875 ,n930);
    or g1266(n1386 ,n1119 ,n1192);
    or g1267(n1385 ,n1183 ,n1182);
    or g1268(n1384 ,n1179 ,n1178);
    or g1269(n1383 ,n653 ,n1189);
    or g1270(n1382 ,n1180 ,n1177);
    or g1271(n1381 ,n782 ,n1076);
    or g1272(n1380 ,n1176 ,n1174);
    or g1273(n1379 ,n680 ,n905);
    or g1274(n1378 ,n677 ,n906);
    or g1275(n1377 ,n676 ,n907);
    or g1276(n1376 ,n1171 ,n1170);
    or g1277(n1375 ,n678 ,n908);
    or g1278(n1374 ,n674 ,n909);
    or g1279(n1373 ,n679 ,n910);
    or g1280(n1372 ,n675 ,n784);
    or g1281(n1371 ,n896 ,n947);
    or g1282(n1370 ,n652 ,n1166);
    or g1283(n1369 ,n1165 ,n1164);
    or g1284(n1368 ,n858 ,n931);
    or g1285(n1367 ,n655 ,n1194);
    or g1286(n1366 ,n857 ,n1060);
    or g1287(n1365 ,n870 ,n1059);
    or g1288(n1364 ,n1163 ,n1162);
    or g1289(n1363 ,n877 ,n1057);
    or g1290(n1362 ,n862 ,n952);
    or g1291(n1361 ,n879 ,n1056);
    or g1292(n1360 ,n854 ,n1055);
    or g1293(n1359 ,n884 ,n1054);
    or g1294(n1358 ,n1209 ,n1196);
    or g1295(n1357 ,n853 ,n1053);
    or g1296(n1356 ,n1159 ,n1158);
    or g1297(n1355 ,n849 ,n1051);
    or g1298(n1354 ,n893 ,n1049);
    or g1299(n1353 ,n787 ,n1048);
    or g1300(n1352 ,n848 ,n1047);
    or g1301(n1351 ,n898 ,n1046);
    or g1302(n1350 ,n847 ,n1045);
    or g1303(n1349 ,n904 ,n1044);
    or g1304(n1348 ,n1157 ,n1156);
    or g1305(n1347 ,n1155 ,n1154);
    or g1306(n1346 ,n812 ,n1042);
    or g1307(n1345 ,n843 ,n1041);
    or g1308(n1344 ,n1167 ,n1204);
    or g1309(n1343 ,n864 ,n1065);
    or g1310(n1342 ,n1152 ,n1151);
    or g1311(n1341 ,n842 ,n1040);
    or g1312(n1340 ,n841 ,n1039);
    or g1313(n1339 ,n840 ,n1038);
    or g1314(n1338 ,n883 ,n1037);
    or g1315(n1337 ,n837 ,n1035);
    or g1316(n1336 ,n894 ,n1034);
    or g1317(n1335 ,n836 ,n1073);
    or g1318(n1334 ,n897 ,n1033);
    or g1319(n1333 ,n801 ,n1031);
    or g1320(n1332 ,n892 ,n1030);
    or g1321(n1331 ,n835 ,n1029);
    or g1322(n1330 ,n650 ,n1148);
    or g1323(n1329 ,n1147 ,n1146);
    or g1324(n1328 ,n832 ,n1026);
    or g1325(n1327 ,n796 ,n942);
    or g1326(n1326 ,n790 ,n1024);
    or g1327(n1325 ,n1145 ,n1143);
    or g1328(n1324 ,n831 ,n1023);
    or g1329(n1323 ,n830 ,n1022);
    or g1330(n1322 ,n800 ,n1021);
    or g1331(n1321 ,n829 ,n1020);
    or g1332(n1320 ,n1207 ,n1130);
    or g1333(n1319 ,n872 ,n932);
    or g1334(n1318 ,n827 ,n1018);
    or g1335(n1317 ,n865 ,n1066);
    or g1336(n1316 ,n860 ,n1028);
    or g1337(n1315 ,n826 ,n1017);
    or g1338(n1314 ,n895 ,n1016);
    or g1339(n1313 ,n1140 ,n1139);
    or g1340(n1312 ,n825 ,n1015);
    or g1341(n1311 ,n863 ,n1068);
    or g1342(n1310 ,n871 ,n1012);
    or g1343(n1309 ,n789 ,n1010);
    or g1344(n1308 ,n1137 ,n1136);
    or g1345(n1307 ,n822 ,n1009);
    or g1346(n1306 ,n833 ,n1008);
    or g1347(n1305 ,n819 ,n940);
    or g1348(n1304 ,n816 ,n1007);
    or g1349(n1303 ,n1133 ,n1132);
    or g1350(n1302 ,n903 ,n1006);
    or g1351(n1301 ,n861 ,n1005);
    or g1352(n1300 ,n811 ,n936);
    or g1353(n1299 ,n1131 ,n1129);
    or g1354(n1298 ,n873 ,n957);
    or g1355(n1297 ,n802 ,n1226);
    or g1356(n1296 ,n815 ,n976);
    or g1357(n1295 ,n886 ,n974);
    or g1358(n1294 ,n651 ,n1124);
    or g1359(n1293 ,n882 ,n973);
    or g1360(n1292 ,n1213 ,n1211);
    or g1361(n1291 ,n902 ,n972);
    or g1362(n1290 ,n869 ,n970);
    or g1363(n1289 ,n1118 ,n1112);
    or g1364(n1288 ,n785 ,n968);
    or g1365(n1287 ,n649 ,n1123);
    or g1366(n1286 ,n810 ,n967);
    or g1367(n1285 ,n1121 ,n1120);
    or g1368(n1284 ,n791 ,n966);
    or g1369(n1283 ,n803 ,n945);
    or g1370(n1282 ,n792 ,n965);
    or g1371(n1281 ,n794 ,n964);
    or g1372(n1280 ,n808 ,n963);
    or g1373(n1279 ,n1127 ,n1134);
    or g1374(n1278 ,n799 ,n962);
    or g1375(n1277 ,n1116 ,n1227);
    or g1376(n1276 ,n821 ,n960);
    or g1377(n1275 ,n813 ,n971);
    or g1378(n1274 ,n817 ,n959);
    or g1379(n1273 ,n820 ,n958);
    or g1380(n1272 ,n805 ,n1013);
    or g1381(n1271 ,n818 ,n969);
    or g1382(n1270 ,n683 ,n1220);
    or g1383(n1269 ,n900 ,n956);
    or g1384(n1268 ,n1109 ,n1110);
    or g1385(n1267 ,n850 ,n954);
    or g1386(n1266 ,n852 ,n1050);
    or g1387(n1265 ,n1168 ,n1108);
    or g1388(n1264 ,n855 ,n953);
    or g1389(n1263 ,n846 ,n937);
    or g1390(n1262 ,n804 ,n951);
    or g1391(n1261 ,n899 ,n1075);
    or g1392(n1260 ,n1106 ,n1105);
    or g1393(n1259 ,n1107 ,n1100);
    or g1394(n1258 ,n1102 ,n1113);
    or g1395(n1257 ,n890 ,n949);
    or g1396(n1256 ,n1103 ,n1101);
    or g1397(n1255 ,n806 ,n948);
    or g1398(n1254 ,n657 ,n1128);
    or g1399(n1253 ,n867 ,n946);
    or g1400(n1252 ,n795 ,n1063);
    or g1401(n1251 ,n881 ,n1067);
    or g1402(n1250 ,n1093 ,n1111);
    or g1403(n1249 ,n888 ,n944);
    or g1404(n1248 ,n891 ,n943);
    or g1405(n1247 ,n885 ,n1064);
    or g1406(n1246 ,n874 ,n941);
    or g1407(n1245 ,n786 ,n939);
    or g1408(n1244 ,n788 ,n938);
    or g1409(n1243 ,n656 ,n1098);
    or g1410(n1242 ,n793 ,n934);
    or g1411(n1241 ,n1097 ,n1096);
    or g1412(n1240 ,n732 ,n1225);
    or g1413(n1239 ,n809 ,n935);
    or g1414(n1238 ,n814 ,n975);
    or g1415(n1237 ,n824 ,n933);
    or g1416(n1236 ,n1138 ,n1188);
    or g1417(n1235 ,n1095 ,n1092);
    or g1418(n1234 ,n844 ,n925);
    or g1419(n1233 ,n1089 ,n1212);
    or g1420(n1232 ,n856 ,n1058);
    or g1421(n1231 ,n1200 ,n1206);
    or g1422(n1230 ,n880 ,n1069);
    or g1423(n1229 ,n889 ,n929);
    or g1424(n1228 ,n1088 ,n1191);
    nor g1425(n1412 ,n517 ,n996);
    nor g1426(n1410 ,n586 ,n996);
    nor g1427(n1227 ,n193 ,n770);
    nor g1428(n1226 ,n250 ,n691);
    nor g1429(n1225 ,n170 ,n717);
    nor g1430(n1224 ,n343 ,n718);
    nor g1431(n1223 ,n346 ,n717);
    nor g1432(n1222 ,n350 ,n717);
    nor g1433(n1221 ,n340 ,n718);
    nor g1434(n1220 ,n168 ,n717);
    nor g1435(n1219 ,n351 ,n716);
    nor g1436(n1218 ,n349 ,n716);
    nor g1437(n1217 ,n344 ,n716);
    nor g1438(n1216 ,n348 ,n716);
    nor g1439(n1215 ,n275 ,n767);
    nor g1440(n1214 ,n239 ,n752);
    nor g1441(n1213 ,n356 ,n767);
    nor g1442(n1212 ,n195 ,n689);
    nor g1443(n1211 ,n437 ,n761);
    nor g1444(n1210 ,n456 ,n709);
    nor g1445(n1209 ,n400 ,n754);
    nor g1446(n1208 ,n200 ,n709);
    nor g1447(n1207 ,n477 ,n758);
    nor g1448(n1206 ,n406 ,n769);
    nor g1449(n1205 ,n270 ,n770);
    nor g1450(n1204 ,n374 ,n770);
    nor g1451(n1203 ,n368 ,n759);
    nor g1452(n1202 ,n291 ,n709);
    nor g1453(n1201 ,n254 ,n769);
    nor g1454(n1200 ,n466 ,n698);
    nor g1455(n1199 ,n187 ,n709);
    nor g1456(n1198 ,n465 ,n751);
    nor g1457(n1197 ,n402 ,n758);
    nor g1458(n1196 ,n185 ,n752);
    nor g1459(n1195 ,n436 ,n758);
    nor g1460(n1194 ,n244 ,n713);
    nor g1461(n1193 ,n279 ,n709);
    nor g1462(n1192 ,n260 ,n689);
    nor g1463(n1191 ,n202 ,n689);
    nor g1464(n1190 ,n204 ,n698);
    nor g1465(n1189 ,n354 ,n713);
    nor g1466(n1188 ,n175 ,n769);
    nor g1467(n1187 ,n214 ,n706);
    nor g1468(n1186 ,n385 ,n709);
    nor g1469(n1185 ,n295 ,n706);
    nor g1470(n1184 ,n221 ,n751);
    nor g1471(n1183 ,n183 ,n767);
    nor g1472(n1182 ,n230 ,n761);
    nor g1473(n1181 ,n268 ,n769);
    nor g1474(n1180 ,n236 ,n754);
    nor g1475(n1179 ,n424 ,n749);
    nor g1476(n1178 ,n438 ,n689);
    nor g1477(n1177 ,n416 ,n752);
    nor g1478(n1176 ,n381 ,n767);
    nor g1479(n1175 ,n358 ,n698);
    nor g1480(n1174 ,n371 ,n761);
    nor g1481(n1173 ,n232 ,n769);
    nor g1482(n1172 ,n510 ,n751);
    nor g1483(n1171 ,n393 ,n754);
    nor g1484(n1170 ,n479 ,n752);
    nor g1485(n1169 ,n501 ,n751);
    nor g1486(n1168 ,n418 ,n749);
    nor g1487(n1167 ,n205 ,n753);
    nor g1488(n1166 ,n447 ,n713);
    nor g1489(n1165 ,n282 ,n758);
    nor g1490(n1164 ,n484 ,n759);
    nor g1491(n1163 ,n495 ,n753);
    nor g1492(n1162 ,n219 ,n770);
    nor g1493(n1161 ,n247 ,n706);
    nor g1494(n1160 ,n488 ,n706);
    nor g1495(n1159 ,n467 ,n698);
    nor g1496(n1158 ,n257 ,n769);
    nor g1497(n1157 ,n398 ,n749);
    nor g1498(n1156 ,n425 ,n689);
    nor g1499(n1155 ,n287 ,n767);
    nor g1500(n1154 ,n417 ,n761);
    nor g1501(n1153 ,n365 ,n751);
    nor g1502(n1152 ,n357 ,n754);
    nor g1503(n1151 ,n208 ,n752);
    nor g1504(n1150 ,n459 ,n751);
    nor g1505(n1149 ,n176 ,n753);
    nor g1506(n1148 ,n382 ,n713);
    nor g1507(n1147 ,n182 ,n758);
    nor g1508(n1146 ,n281 ,n759);
    nor g1509(n1145 ,n474 ,n753);
    nor g1510(n1144 ,n396 ,n770);
    nor g1511(n1143 ,n363 ,n770);
    nor g1512(n1142 ,n197 ,n751);
    nor g1513(n1141 ,n475 ,n706);
    nor g1514(n1140 ,n509 ,n698);
    nor g1515(n1139 ,n217 ,n769);
    nor g1516(n1138 ,n497 ,n698);
    nor g1517(n1137 ,n485 ,n749);
    nor g1518(n1136 ,n405 ,n689);
    nor g1519(n1135 ,n428 ,n698);
    nor g1520(n1134 ,n234 ,n752);
    nor g1521(n1133 ,n472 ,n767);
    nor g1522(n1132 ,n361 ,n761);
    nor g1523(n1131 ,n390 ,n754);
    nor g1524(n1130 ,n194 ,n759);
    nor g1525(n1129 ,n468 ,n752);
    nor g1526(n1128 ,n226 ,n713);
    nor g1527(n1127 ,n434 ,n754);
    nor g1528(n1126 ,n243 ,n751);
    nor g1529(n1125 ,n409 ,n709);
    nor g1530(n1124 ,n464 ,n713);
    nor g1531(n1123 ,n470 ,n713);
    nor g1532(n1122 ,n375 ,n709);
    nor g1533(n1121 ,n491 ,n758);
    nor g1534(n1120 ,n276 ,n759);
    nor g1535(n1119 ,n442 ,n749);
    nor g1536(n1118 ,n432 ,n758);
    nor g1537(n1117 ,n177 ,n759);
    nor g1538(n1116 ,n191 ,n753);
    nor g1539(n1115 ,n256 ,n691);
    nor g1540(n1114 ,n391 ,n706);
    nor g1541(n1113 ,n384 ,n761);
    nor g1542(n1112 ,n503 ,n759);
    nor g1543(n1111 ,n461 ,n689);
    nor g1544(n1110 ,n378 ,n769);
    nor g1545(n1109 ,n455 ,n698);
    nor g1546(n1108 ,n430 ,n689);
    nor g1547(n1107 ,n476 ,n753);
    nor g1548(n1106 ,n292 ,n767);
    nor g1549(n1105 ,n453 ,n761);
    nor g1550(n1104 ,n389 ,n754);
    nor g1551(n1103 ,n245 ,n754);
    nor g1552(n1102 ,n370 ,n767);
    nor g1553(n1101 ,n421 ,n752);
    nor g1554(n1100 ,n273 ,n770);
    nor g1555(n1099 ,n284 ,n753);
    nor g1556(n1098 ,n478 ,n713);
    nor g1557(n1097 ,n209 ,n758);
    nor g1558(n1096 ,n469 ,n759);
    nor g1559(n1095 ,n203 ,n753);
    nor g1560(n1094 ,n379 ,n706);
    nor g1561(n1093 ,n222 ,n749);
    nor g1562(n1092 ,n502 ,n770);
    nor g1563(n1091 ,n408 ,n761);
    nor g1564(n1090 ,n395 ,n706);
    nor g1565(n1089 ,n251 ,n749);
    nor g1566(n1088 ,n493 ,n749);
    nor g1567(n1087 ,n376 ,n748);
    nor g1568(n1086 ,n360 ,n748);
    nor g1569(n1085 ,n494 ,n748);
    nor g1570(n1084 ,n218 ,n748);
    nor g1571(n1083 ,n355 ,n748);
    nor g1572(n1082 ,n407 ,n748);
    nor g1573(n1081 ,n367 ,n748);
    nor g1574(n1080 ,n399 ,n748);
    nor g1575(n1079 ,n392 ,n711);
    nor g1576(n1078 ,n179 ,n711);
    nor g1577(n1077 ,n420 ,n711);
    nor g1578(n1076 ,n440 ,n711);
    nor g1579(n1075 ,n252 ,n697);
    nor g1580(n1074 ,n482 ,n693);
    nor g1581(n1073 ,n489 ,n703);
    nor g1582(n1072 ,n435 ,n707);
    nor g1583(n1071 ,n269 ,n690);
    nor g1584(n1070 ,n415 ,n708);
    nor g1585(n1069 ,n496 ,n690);
    nor g1586(n1068 ,n404 ,n694);
    nor g1587(n1067 ,n504 ,n692);
    nor g1588(n1066 ,n401 ,n694);
    nor g1589(n1065 ,n294 ,n700);
    nor g1590(n1064 ,n290 ,n708);
    nor g1591(n1063 ,n383 ,n692);
    nor g1592(n1062 ,n500 ,n692);
    nor g1593(n1061 ,n450 ,n702);
    nor g1594(n1060 ,n283 ,n702);
    nor g1595(n1059 ,n353 ,n702);
    nor g1596(n1058 ,n253 ,n690);
    nor g1597(n1057 ,n481 ,n702);
    nor g1598(n1056 ,n241 ,n702);
    nor g1599(n1055 ,n263 ,n702);
    nor g1600(n1054 ,n366 ,n702);
    nor g1601(n1053 ,n249 ,n702);
    nor g1602(n1052 ,n190 ,n701);
    nor g1603(n1051 ,n498 ,n701);
    nor g1604(n1050 ,n231 ,n697);
    nor g1605(n1049 ,n506 ,n701);
    nor g1606(n1048 ,n278 ,n701);
    nor g1607(n1047 ,n423 ,n701);
    nor g1608(n1046 ,n215 ,n701);
    nor g1609(n1045 ,n422 ,n701);
    nor g1610(n1044 ,n487 ,n701);
    nor g1611(n1043 ,n471 ,n700);
    nor g1612(n1042 ,n277 ,n700);
    nor g1613(n1041 ,n448 ,n700);
    nor g1614(n1040 ,n206 ,n700);
    nor g1615(n1039 ,n433 ,n700);
    nor g1616(n1038 ,n271 ,n700);
    nor g1617(n1037 ,n446 ,n700);
    nor g1618(n1036 ,n499 ,n703);
    nor g1619(n1035 ,n262 ,n703);
    nor g1620(n1034 ,n380 ,n703);
    nor g1621(n1033 ,n439 ,n703);
    nor g1622(n1032 ,n431 ,n690);
    nor g1623(n1031 ,n457 ,n703);
    nor g1624(n1030 ,n228 ,n703);
    nor g1625(n1029 ,n373 ,n703);
    nor g1626(n1028 ,n445 ,n707);
    nor g1627(n1027 ,n288 ,n696);
    nor g1628(n1026 ,n427 ,n696);
    nor g1629(n1025 ,n180 ,n711);
    nor g1630(n1024 ,n267 ,n696);
    nor g1631(n1023 ,n285 ,n696);
    nor g1632(n1022 ,n213 ,n696);
    nor g1633(n1021 ,n181 ,n696);
    nor g1634(n1020 ,n255 ,n696);
    nor g1635(n1019 ,n352 ,n694);
    nor g1636(n1018 ,n274 ,n694);
    nor g1637(n1017 ,n237 ,n694);
    nor g1638(n1016 ,n233 ,n694);
    nor g1639(n1015 ,n452 ,n694);
    nor g1640(n1014 ,n369 ,n711);
    nor g1641(n1013 ,n443 ,n695);
    nor g1642(n1012 ,n410 ,n694);
    nor g1643(n1011 ,n266 ,n710);
    nor g1644(n1010 ,n186 ,n710);
    nor g1645(n1009 ,n429 ,n710);
    nor g1646(n1008 ,n480 ,n710);
    nor g1647(n1007 ,n412 ,n710);
    nor g1648(n1006 ,n261 ,n710);
    nor g1649(n1005 ,n289 ,n710);
    not g1650(n1003 ,n1002);
    not g1651(n995 ,n996);
    not g1652(n979 ,n978);
    or g1653(n977 ,n660 ,n735);
    nor g1654(n976 ,n508 ,n691);
    nor g1655(n975 ,n272 ,n707);
    nor g1656(n974 ,n507 ,n691);
    nor g1657(n973 ,n265 ,n691);
    nor g1658(n972 ,n463 ,n691);
    nor g1659(n971 ,n426 ,n695);
    nor g1660(n970 ,n413 ,n691);
    nor g1661(n969 ,n386 ,n695);
    nor g1662(n968 ,n199 ,n693);
    nor g1663(n967 ,n394 ,n693);
    nor g1664(n966 ,n238 ,n693);
    nor g1665(n965 ,n258 ,n693);
    nor g1666(n964 ,n490 ,n693);
    nor g1667(n963 ,n264 ,n693);
    nor g1668(n962 ,n259 ,n693);
    nor g1669(n961 ,n212 ,n695);
    nor g1670(n960 ,n454 ,n695);
    nor g1671(n959 ,n201 ,n695);
    nor g1672(n958 ,n240 ,n695);
    nor g1673(n957 ,n505 ,n691);
    nor g1674(n956 ,n280 ,n695);
    nor g1675(n955 ,n483 ,n697);
    nor g1676(n954 ,n286 ,n697);
    nor g1677(n953 ,n473 ,n697);
    nor g1678(n952 ,n414 ,n697);
    nor g1679(n951 ,n248 ,n697);
    nor g1680(n950 ,n449 ,n697);
    nor g1681(n949 ,n364 ,n692);
    nor g1682(n948 ,n362 ,n692);
    nor g1683(n947 ,n293 ,n692);
    nor g1684(n946 ,n397 ,n692);
    nor g1685(n945 ,n387 ,n692);
    nor g1686(n944 ,n359 ,n708);
    nor g1687(n943 ,n224 ,n708);
    nor g1688(n942 ,n372 ,n696);
    nor g1689(n941 ,n210 ,n708);
    nor g1690(n940 ,n492 ,n710);
    nor g1691(n939 ,n486 ,n708);
    nor g1692(n938 ,n207 ,n708);
    nor g1693(n937 ,n220 ,n707);
    nor g1694(n936 ,n184 ,n707);
    nor g1695(n935 ,n419 ,n707);
    nor g1696(n934 ,n174 ,n708);
    nor g1697(n933 ,n377 ,n707);
    nor g1698(n932 ,n411 ,n707);
    nor g1699(n931 ,n444 ,n690);
    nor g1700(n930 ,n225 ,n690);
    nor g1701(n929 ,n246 ,n690);
    nor g1702(n928 ,n223 ,n711);
    nor g1703(n927 ,n458 ,n711);
    nor g1704(n926 ,n338 ,n718);
    nor g1705(n925 ,n242 ,n690);
    or g1706(n924 ,n563 ,n724);
    nor g1707(n923 ,n330 ,n718);
    nor g1708(n922 ,n162 ,n716);
    or g1709(n921 ,n641 ,n729);
    or g1710(n920 ,n658 ,n733);
    or g1711(n919 ,n662 ,n734);
    or g1712(n918 ,n659 ,n736);
    nor g1713(n917 ,n142 ,n686);
    nor g1714(n916 ,n142 ,n687);
    nor g1715(n915 ,n527 ,n715);
    or g1716(n914 ,n579 ,n682);
    or g1717(n913 ,n585 ,n681);
    or g1718(n912 ,n578 ,n672);
    or g1719(n911 ,n577 ,n673);
    nor g1720(n910 ,n150 ,n714);
    nor g1721(n909 ,n329 ,n714);
    nor g1722(n908 ,n327 ,n714);
    nor g1723(n907 ,n328 ,n714);
    nor g1724(n906 ,n148 ,n714);
    nor g1725(n905 ,n149 ,n714);
    nor g1726(n904 ,n154 ,n765);
    nor g1727(n903 ,n156 ,n704);
    nor g1728(n902 ,n156 ,n750);
    nor g1729(n901 ,n154 ,n764);
    nor g1730(n900 ,n154 ,n699);
    nor g1731(n899 ,n156 ,n764);
    nor g1732(n898 ,n157 ,n765);
    nor g1733(n897 ,n153 ,n768);
    nor g1734(n896 ,n155 ,n760);
    nor g1735(n895 ,n153 ,n712);
    nor g1736(n894 ,n158 ,n768);
    nor g1737(n893 ,n158 ,n765);
    nor g1738(n892 ,n156 ,n768);
    nor g1739(n891 ,n158 ,n763);
    nor g1740(n890 ,n159 ,n760);
    nor g1741(n889 ,n154 ,n755);
    nor g1742(n888 ,n159 ,n763);
    nor g1743(n887 ,n156 ,n755);
    nor g1744(n886 ,n153 ,n750);
    nor g1745(n885 ,n155 ,n763);
    nor g1746(n884 ,n156 ,n757);
    nor g1747(n883 ,n154 ,n756);
    nor g1748(n882 ,n157 ,n750);
    nor g1749(n881 ,n154 ,n760);
    nor g1750(n880 ,n157 ,n755);
    nor g1751(n879 ,n153 ,n757);
    nor g1752(n878 ,n152 ,n764);
    nor g1753(n877 ,n155 ,n757);
    nor g1754(n876 ,n152 ,n763);
    nor g1755(n875 ,n153 ,n755);
    nor g1756(n874 ,n153 ,n763);
    nor g1757(n873 ,n159 ,n750);
    nor g1758(n872 ,n154 ,n766);
    nor g1759(n871 ,n154 ,n712);
    nor g1760(n870 ,n158 ,n757);
    nor g1761(n869 ,n154 ,n750);
    nor g1762(n868 ,n152 ,n750);
    nor g1763(n867 ,n153 ,n760);
    nor g1764(n866 ,n152 ,n762);
    nor g1765(n865 ,n158 ,n712);
    nor g1766(n864 ,n155 ,n756);
    nor g1767(n863 ,n156 ,n712);
    nor g1768(n862 ,n153 ,n764);
    nor g1769(n861 ,n154 ,n704);
    nor g1770(n860 ,n156 ,n766);
    nor g1771(n859 ,n152 ,n757);
    nor g1772(n858 ,n155 ,n755);
    nor g1773(n857 ,n159 ,n757);
    nor g1774(n856 ,n158 ,n755);
    nor g1775(n855 ,n155 ,n764);
    nor g1776(n854 ,n157 ,n757);
    nor g1777(n853 ,n154 ,n757);
    nor g1778(n852 ,n158 ,n764);
    nor g1779(n851 ,n152 ,n765);
    nor g1780(n850 ,n159 ,n764);
    nor g1781(n849 ,n159 ,n765);
    nor g1782(n848 ,n153 ,n765);
    nor g1783(n847 ,n156 ,n765);
    nor g1784(n846 ,n159 ,n766);
    nor g1785(n845 ,n152 ,n756);
    nor g1786(n844 ,n159 ,n755);
    nor g1787(n843 ,n158 ,n756);
    nor g1788(n842 ,n153 ,n756);
    nor g1789(n841 ,n157 ,n756);
    nor g1790(n840 ,n156 ,n756);
    nor g1791(n839 ,n152 ,n755);
    nor g1792(n838 ,n152 ,n768);
    nor g1793(n837 ,n159 ,n768);
    nor g1794(n836 ,n155 ,n768);
    nor g1795(n835 ,n154 ,n768);
    nor g1796(n834 ,n152 ,n705);
    nor g1797(n833 ,n155 ,n704);
    nor g1798(n832 ,n159 ,n705);
    nor g1799(n831 ,n153 ,n705);
    nor g1800(n830 ,n157 ,n705);
    nor g1801(n829 ,n154 ,n705);
    nor g1802(n828 ,n152 ,n712);
    nor g1803(n827 ,n159 ,n712);
    nor g1804(n826 ,n155 ,n712);
    nor g1805(n825 ,n157 ,n712);
    nor g1806(n824 ,n157 ,n766);
    nor g1807(n823 ,n152 ,n704);
    nor g1808(n822 ,n158 ,n704);
    nor g1809(n821 ,n159 ,n699);
    nor g1810(n820 ,n153 ,n699);
    nor g1811(n819 ,n153 ,n704);
    nor g1812(n818 ,n156 ,n699);
    nor g1813(n817 ,n155 ,n699);
    nor g1814(n816 ,n157 ,n704);
    nor g1815(n815 ,n155 ,n750);
    nor g1816(n814 ,n153 ,n766);
    nor g1817(n813 ,n158 ,n699);
    nor g1818(n812 ,n159 ,n756);
    nor g1819(n811 ,n158 ,n766);
    nor g1820(n810 ,n158 ,n762);
    nor g1821(n809 ,n155 ,n766);
    nor g1822(n808 ,n156 ,n762);
    nor g1823(n807 ,n152 ,n699);
    nor g1824(n806 ,n158 ,n760);
    nor g1825(n805 ,n157 ,n699);
    nor g1826(n804 ,n157 ,n764);
    nor g1827(n803 ,n157 ,n760);
    nor g1828(n802 ,n158 ,n750);
    nor g1829(n801 ,n157 ,n768);
    nor g1830(n800 ,n156 ,n705);
    nor g1831(n799 ,n154 ,n762);
    nor g1832(n798 ,n152 ,n760);
    nor g1833(n797 ,n152 ,n766);
    nor g1834(n796 ,n158 ,n705);
    nor g1835(n795 ,n156 ,n760);
    nor g1836(n794 ,n157 ,n762);
    nor g1837(n793 ,n154 ,n763);
    nor g1838(n792 ,n153 ,n762);
    nor g1839(n791 ,n155 ,n762);
    nor g1840(n790 ,n155 ,n705);
    nor g1841(n789 ,n159 ,n704);
    nor g1842(n788 ,n156 ,n763);
    nor g1843(n787 ,n155 ,n765);
    nor g1844(n786 ,n157 ,n763);
    nor g1845(n785 ,n159 ,n762);
    nor g1846(n784 ,n151 ,n714);
    nor g1847(n783 ,n154 ,n746);
    nor g1848(n782 ,n159 ,n746);
    nor g1849(n781 ,n158 ,n746);
    nor g1850(n780 ,n156 ,n746);
    nor g1851(n779 ,n157 ,n746);
    nor g1852(n778 ,n153 ,n746);
    nor g1853(n777 ,n155 ,n746);
    nor g1854(n776 ,n152 ,n746);
    nor g1855(n1002 ,n643 ,n725);
    or g1856(n1001 ,n626 ,n745);
    or g1857(n1000 ,n334 ,n723);
    or g1858(n999 ,n38[2] ,n723);
    or g1859(n998 ,n38[2] ,n775);
    or g1860(n997 ,n334 ,n775);
    nor g1861(n996 ,n36[4] ,n726);
    or g1862(n994 ,n520 ,n774);
    or g1863(n993 ,n534 ,n722);
    or g1864(n992 ,n538 ,n721);
    or g1865(n991 ,n520 ,n722);
    or g1866(n990 ,n522 ,n722);
    or g1867(n989 ,n538 ,n774);
    or g1868(n988 ,n534 ,n721);
    or g1869(n987 ,n534 ,n772);
    or g1870(n986 ,n534 ,n774);
    or g1871(n985 ,n520 ,n772);
    or g1872(n984 ,n522 ,n772);
    or g1873(n983 ,n522 ,n721);
    or g1874(n982 ,n538 ,n722);
    or g1875(n981 ,n520 ,n721);
    or g1876(n980 ,n522 ,n774);
    nor g1877(n978 ,n538 ,n772);
    not g1878(n748 ,n747);
    not g1879(n746 ,n745);
    nor g1880(n744 ,n164 ,n629);
    nor g1881(n743 ,n409 ,n628);
    nor g1882(n742 ,n291 ,n628);
    nor g1883(n741 ,n375 ,n628);
    nor g1884(n740 ,n279 ,n628);
    nor g1885(n739 ,n200 ,n628);
    nor g1886(n738 ,n385 ,n628);
    nor g1887(n737 ,n456 ,n628);
    nor g1888(n736 ,n303 ,n626);
    nor g1889(n735 ,n323 ,n626);
    nor g1890(n734 ,n305 ,n626);
    nor g1891(n733 ,n298 ,n626);
    nor g1892(n732 ,n315 ,n624);
    nor g1893(n731 ,n299 ,n624);
    nor g1894(n730 ,n316 ,n624);
    nor g1895(n729 ,n341 ,n629);
    nor g1896(n728 ,n333 ,n629);
    nor g1897(n727 ,n336 ,n629);
    or g1898(n775 ,n342 ,n647);
    or g1899(n774 ,n336 ,n642);
    or g1900(n773 ,n166 ,n646);
    or g1901(n772 ,n336 ,n670);
    or g1902(n771 ,n166 ,n671);
    or g1903(n770 ,n535 ,n669);
    or g1904(n769 ,n523 ,n669);
    or g1905(n768 ,n559 ,n637);
    or g1906(n767 ,n537 ,n638);
    or g1907(n766 ,n572 ,n635);
    or g1908(n765 ,n559 ,n640);
    or g1909(n764 ,n558 ,n636);
    or g1910(n763 ,n571 ,n635);
    or g1911(n762 ,n558 ,n635);
    or g1912(n761 ,n537 ,n639);
    or g1913(n760 ,n559 ,n636);
    or g1914(n759 ,n537 ,n669);
    or g1915(n758 ,n537 ,n668);
    or g1916(n757 ,n558 ,n640);
    or g1917(n756 ,n558 ,n637);
    or g1918(n755 ,n571 ,n636);
    or g1919(n754 ,n523 ,n638);
    or g1920(n753 ,n535 ,n668);
    or g1921(n752 ,n523 ,n639);
    or g1922(n751 ,n523 ,n668);
    or g1923(n750 ,n572 ,n637);
    or g1924(n749 ,n535 ,n638);
    nor g1925(n747 ,n539 ,n668);
    nor g1926(n745 ,n572 ,n636);
    not g1927(n725 ,n724);
    not g1928(n716 ,n715);
    nor g1929(n688 ,n59[0] ,n626);
    nor g1930(n687 ,n663 ,n620);
    nor g1931(n686 ,n648 ,n664);
    or g1932(n685 ,n625 ,n654);
    or g1933(n684 ,n592 ,n667);
    nor g1934(n683 ,n18[0] ,n624);
    or g1935(n682 ,n568 ,n631);
    or g1936(n681 ,n565 ,n631);
    nor g1937(n680 ,n2296 ,n624);
    nor g1938(n679 ,n329 ,n624);
    nor g1939(n678 ,n328 ,n624);
    nor g1940(n677 ,n149 ,n624);
    nor g1941(n676 ,n148 ,n624);
    nor g1942(n675 ,n150 ,n624);
    nor g1943(n674 ,n327 ,n624);
    or g1944(n673 ,n567 ,n631);
    or g1945(n672 ,n566 ,n631);
    or g1946(n726 ,n15 ,n645);
    nor g1947(n724 ,n564 ,n644);
    or g1948(n723 ,n38[1] ,n647);
    or g1949(n722 ,n58[3] ,n642);
    or g1950(n721 ,n58[3] ,n670);
    or g1951(n720 ,n38[3] ,n646);
    or g1952(n719 ,n38[3] ,n671);
    or g1953(n718 ,n145 ,n627);
    or g1954(n717 ,n557 ,n625);
    nor g1955(n715 ,n627 ,n629);
    or g1956(n714 ,n145 ,n625);
    or g1957(n713 ,n539 ,n638);
    or g1958(n712 ,n572 ,n640);
    nor g1959(n711 ,n633 ,n591);
    nor g1960(n710 ,n633 ,n588);
    or g1961(n709 ,n611 ,n629);
    nor g1962(n708 ,n634 ,n590);
    nor g1963(n707 ,n591 ,n634);
    or g1964(n706 ,n539 ,n669);
    or g1965(n705 ,n571 ,n640);
    or g1966(n704 ,n571 ,n637);
    nor g1967(n703 ,n630 ,n589);
    nor g1968(n702 ,n632 ,n588);
    nor g1969(n701 ,n589 ,n632);
    nor g1970(n700 ,n630 ,n588);
    or g1971(n699 ,n559 ,n635);
    or g1972(n698 ,n539 ,n639);
    nor g1973(n697 ,n630 ,n590);
    nor g1974(n696 ,n634 ,n588);
    nor g1975(n695 ,n591 ,n632);
    nor g1976(n694 ,n634 ,n589);
    nor g1977(n693 ,n590 ,n632);
    nor g1978(n692 ,n591 ,n630);
    nor g1979(n691 ,n633 ,n589);
    nor g1980(n690 ,n633 ,n590);
    or g1981(n689 ,n535 ,n639);
    nor g1982(n667 ,n167 ,n586);
    nor g1983(n666 ,n162 ,n613);
    nor g1984(n665 ,n2297 ,n580);
    nor g1985(n664 ,n187 ,n612);
    nor g1986(n663 ,n462 ,n595);
    nor g1987(n662 ,n306 ,n587);
    nor g1988(n661 ,n163 ,n617);
    nor g1989(n660 ,n324 ,n587);
    nor g1990(n659 ,n300 ,n587);
    nor g1991(n658 ,n312 ,n587);
    nor g1992(n657 ,n189 ,n586);
    nor g1993(n656 ,n229 ,n586);
    nor g1994(n655 ,n451 ,n586);
    nor g1995(n654 ,n165 ,n584);
    nor g1996(n653 ,n192 ,n586);
    nor g1997(n652 ,n196 ,n586);
    nor g1998(n651 ,n227 ,n586);
    nor g1999(n650 ,n178 ,n586);
    nor g2000(n649 ,n235 ,n586);
    nor g2001(n648 ,n216 ,n611);
    or g2002(n671 ,n337 ,n614);
    or g2003(n670 ,n341 ,n587);
    or g2004(n669 ,n332 ,n593);
    or g2005(n668 ,n332 ,n601);
    not g2006(n645 ,n644);
    not g2007(n642 ,n641);
    not g2008(n626 ,n627);
    not g2009(n624 ,n625);
    nor g2010(n623 ,n332 ,n586);
    nor g2011(n622 ,n331 ,n586);
    nor g2012(n621 ,n57[4] ,n613);
    nor g2013(n620 ,n541 ,n594);
    nor g2014(n619 ,n36[4] ,n617);
    nor g2015(n618 ,n335 ,n586);
    or g2016(n647 ,n512 ,n600);
    or g2017(n646 ,n38[0] ,n614);
    nor g2018(n644 ,n544 ,n603);
    or g2019(n643 ,n147 ,n602);
    nor g2020(n641 ,n58[0] ,n587);
    or g2021(n640 ,n521 ,n616);
    or g2022(n639 ,n37[3] ,n593);
    or g2023(n638 ,n516 ,n598);
    or g2024(n637 ,n521 ,n615);
    or g2025(n636 ,n540 ,n615);
    or g2026(n635 ,n540 ,n616);
    nor g2027(n634 ,n142 ,n605);
    nor g2028(n633 ,n143 ,n604);
    nor g2029(n632 ,n142 ,n583);
    or g2030(n631 ,n147 ,n595);
    nor g2031(n630 ,n141 ,n582);
    nor g2032(n629 ,n519 ,n596);
    or g2033(n628 ,n144 ,n612);
    nor g2034(n627 ,n142 ,n581);
    nor g2035(n625 ,n142 ,n599);
    not g2036(n612 ,n611);
    nor g2037(n610 ,n318 ,n555);
    nor g2038(n609 ,n319 ,n555);
    nor g2039(n608 ,n296 ,n555);
    nor g2040(n607 ,n317 ,n555);
    nor g2041(n606 ,n19[0] ,n557);
    nor g2042(n605 ,n330 ,n562);
    nor g2043(n604 ,n330 ,n573);
    or g2044(n603 ,n543 ,n561);
    nor g2045(n602 ,n2299 ,n575);
    or g2046(n601 ,n516 ,n574);
    or g2047(n600 ,n146 ,n570);
    or g2048(n599 ,n15 ,n561);
    or g2049(n598 ,n37[3] ,n574);
    or g2050(n617 ,n515 ,n548);
    or g2051(n616 ,n146 ,n562);
    or g2052(n615 ,n146 ,n573);
    or g2053(n614 ,n511 ,n569);
    or g2054(n613 ,n514 ,n547);
    nor g2055(n611 ,n165 ,n561);
    not g2056(n597 ,n596);
    not g2057(n595 ,n594);
    not g2058(n593 ,n592);
    nor g2059(n585 ,n5[2] ,n556);
    or g2060(n584 ,n557 ,n560);
    nor g2061(n583 ,n59[2] ,n562);
    nor g2062(n582 ,n59[2] ,n573);
    or g2063(n581 ,n57[4] ,n575);
    nor g2064(n579 ,n5[3] ,n556);
    nor g2065(n578 ,n5[1] ,n556);
    nor g2066(n577 ,n5[0] ,n556);
    nor g2067(n576 ,n141 ,n553);
    nor g2068(n596 ,n141 ,n564);
    nor g2069(n594 ,n517 ,n563);
    nor g2070(n592 ,n37[0] ,n555);
    nor g2071(n591 ,n141 ,n552);
    nor g2072(n590 ,n142 ,n550);
    nor g2073(n589 ,n143 ,n549);
    nor g2074(n588 ,n143 ,n551);
    or g2075(n587 ,n533 ,n556);
    or g2076(n586 ,n144 ,n554);
    or g2077(n570 ,n339 ,n543);
    or g2078(n569 ,n172 ,n544);
    nor g2079(n568 ,n198 ,n518);
    nor g2080(n567 ,n388 ,n518);
    nor g2081(n566 ,n460 ,n518);
    nor g2082(n565 ,n441 ,n518);
    or g2083(n575 ,n188 ,n516);
    or g2084(n574 ,n167 ,n545);
    or g2085(n573 ,n340 ,n542);
    or g2086(n572 ,n330 ,n536);
    or g2087(n571 ,n330 ,n524);
    not g2088(n561 ,n560);
    not g2089(n555 ,n554);
    nor g2090(n553 ,n531 ,n513);
    nor g2091(n552 ,n536 ,n540);
    nor g2092(n551 ,n524 ,n521);
    nor g2093(n550 ,n540 ,n524);
    nor g2094(n549 ,n536 ,n521);
    or g2095(n548 ,n36[3] ,n529);
    or g2096(n547 ,n57[3] ,n527);
    nor g2097(n564 ,n161 ,n533);
    nor g2098(n563 ,n533 ,n541);
    or g2099(n562 ,n59[1] ,n542);
    nor g2100(n560 ,n533 ,n528);
    or g2101(n559 ,n59[2] ,n536);
    or g2102(n558 ,n59[2] ,n524);
    or g2103(n557 ,n145 ,n517);
    or g2104(n556 ,n40[1] ,n526);
    nor g2105(n554 ,n545 ,n516);
    not g2106(n533 ,n532);
    nor g2107(n531 ,n173 ,n160);
    nor g2108(n530 ,n173 ,n143);
    nor g2109(n546 ,n211 ,n143);
    or g2110(n545 ,n144 ,n2298);
    or g2111(n544 ,n168 ,n350);
    or g2112(n543 ,n170 ,n18[3]);
    or g2113(n542 ,n188 ,n40[0]);
    or g2114(n541 ,n161 ,n160);
    or g2115(n540 ,n343 ,n57[4]);
    or g2116(n539 ,n335 ,n331);
    or g2117(n538 ,n333 ,n164);
    or g2118(n537 ,n335 ,n37[2]);
    or g2119(n536 ,n338 ,n40[1]);
    or g2120(n535 ,n331 ,n37[1]);
    or g2121(n534 ,n164 ,n58[1]);
    nor g2122(n532 ,n339 ,n172);
    not g2123(n526 ,n525);
    not g2124(n518 ,n519);
    not g2125(n516 ,n517);
    or g2126(n515 ,n36[1] ,n36[2]);
    or g2127(n514 ,n57[1] ,n57[2]);
    nor g2128(n513 ,n161 ,n40[1]);
    or g2129(n512 ,n36[4] ,n40[0]);
    or g2130(n511 ,n160 ,n15);
    or g2131(n529 ,n145 ,n36[0]);
    or g2132(n528 ,n160 ,n40[0]);
    or g2133(n527 ,n147 ,n57[0]);
    nor g2134(n525 ,n161 ,n143);
    or g2135(n524 ,n40[1] ,n59[0]);
    or g2136(n523 ,n37[1] ,n37[2]);
    or g2137(n522 ,n58[1] ,n58[2]);
    or g2138(n521 ,n57[4] ,n59[3]);
    or g2139(n520 ,n333 ,n58[2]);
    nor g2140(n519 ,n160 ,n143);
    nor g2141(n517 ,n40[0] ,n40[1]);
    not g2142(n510 ,n29[6]);
    not g2143(n509 ,n26[3]);
    not g2144(n508 ,n48[3]);
    not g2145(n507 ,n48[4]);
    not g2146(n506 ,n42[2]);
    not g2147(n505 ,n48[1]);
    not g2148(n504 ,n52[7]);
    not g2149(n503 ,n30[0]);
    not g2150(n502 ,n32[5]);
    not g2151(n501 ,n29[2]);
    not g2152(n500 ,n52[0]);
    not g2153(n499 ,n44[0]);
    not g2154(n498 ,n42[1]);
    not g2155(n497 ,n26[0]);
    not g2156(n496 ,n55[5]);
    not g2157(n495 ,n33[2]);
    not g2158(n494 ,n35[6]);
    not g2159(n493 ,n25[5]);
    not g2160(n492 ,n47[4]);
    not g2161(n491 ,n31[4]);
    not g2162(n490 ,n49[5]);
    not g2163(n489 ,n44[3]);
    not g2164(n488 ,n34[7]);
    not g2165(n487 ,n42[7]);
    not g2166(n486 ,n53[5]);
    not g2167(n485 ,n25[3]);
    not g2168(n484 ,n30[2]);
    not g2169(n483 ,n51[0]);
    not g2170(n482 ,n49[0]);
    not g2171(n481 ,n41[3]);
    not g2172(n480 ,n47[3]);
    not g2173(n479 ,n20[1]);
    not g2174(n478 ,n27[5]);
    not g2175(n477 ,n31[1]);
    not g2176(n476 ,n33[0]);
    not g2177(n475 ,n34[3]);
    not g2178(n474 ,n33[3]);
    not g2179(n473 ,n51[3]);
    not g2180(n472 ,n23[3]);
    not g2181(n471 ,n43[0]);
    not g2182(n470 ,n27[4]);
    not g2183(n469 ,n30[5]);
    not g2184(n468 ,n20[3]);
    not g2185(n467 ,n26[2]);
    not g2186(n466 ,n26[5]);
    not g2187(n465 ,n29[5]);
    not g2188(n464 ,n27[0]);
    not g2189(n463 ,n48[6]);
    not g2190(n462 ,n11);
    not g2191(n461 ,n24[6]);
    not g2192(n460 ,n17[1]);
    not g2193(n459 ,n29[3]);
    not g2194(n458 ,n56[2]);
    not g2195(n457 ,n44[5]);
    not g2196(n456 ,n60[2]);
    not g2197(n455 ,n26[4]);
    not g2198(n454 ,n50[1]);
    not g2199(n453 ,n22[4]);
    not g2200(n452 ,n46[5]);
    not g2201(n451 ,n6[6]);
    not g2202(n450 ,n41[0]);
    not g2203(n449 ,n51[7]);
    not g2204(n448 ,n43[2]);
    not g2205(n447 ,n27[2]);
    not g2206(n446 ,n43[7]);
    not g2207(n445 ,n54[6]);
    not g2208(n444 ,n55[3]);
    not g2209(n443 ,n50[5]);
    not g2210(n442 ,n25[7]);
    not g2211(n441 ,n17[2]);
    not g2212(n440 ,n56[1]);
    not g2213(n439 ,n44[4]);
    not g2214(n438 ,n24[1]);
    not g2215(n437 ,n22[0]);
    not g2216(n436 ,n31[6]);
    not g2217(n435 ,n54[0]);
    not g2218(n434 ,n21[6]);
    not g2219(n433 ,n43[5]);
    not g2220(n432 ,n31[0]);
    not g2221(n431 ,n55[0]);
    not g2222(n430 ,n24[4]);
    not g2223(n429 ,n47[2]);
    not g2224(n428 ,n26[1]);
    not g2225(n427 ,n45[1]);
    not g2226(n426 ,n50[2]);
    not g2227(n425 ,n24[2]);
    not g2228(n424 ,n25[1]);
    not g2229(n423 ,n42[4]);
    not g2230(n422 ,n42[6]);
    not g2231(n421 ,n20[4]);
    not g2232(n420 ,n56[5]);
    not g2233(n419 ,n54[3]);
    not g2234(n418 ,n25[4]);
    not g2235(n417 ,n22[2]);
    not g2236(n416 ,n20[7]);
    not g2237(n415 ,n53[0]);
    not g2238(n414 ,n51[4]);
    not g2239(n413 ,n48[7]);
    not g2240(n412 ,n47[5]);
    not g2241(n411 ,n54[7]);
    not g2242(n410 ,n46[7]);
    not g2243(n409 ,n60[3]);
    not g2244(n408 ,n22[5]);
    not g2245(n407 ,n35[4]);
    not g2246(n406 ,n28[5]);
    not g2247(n405 ,n24[3]);
    not g2248(n404 ,n46[6]);
    not g2249(n403 ,n12);
    not g2250(n402 ,n31[7]);
    not g2251(n401 ,n46[2]);
    not g2252(n400 ,n21[0]);
    not g2253(n399 ,n35[1]);
    not g2254(n398 ,n25[2]);
    not g2255(n397 ,n52[4]);
    not g2256(n396 ,n32[1]);
    not g2257(n395 ,n34[5]);
    not g2258(n394 ,n49[2]);
    not g2259(n393 ,n21[1]);
    not g2260(n392 ,n56[3]);
    not g2261(n391 ,n34[4]);
    not g2262(n390 ,n21[3]);
    not g2263(n389 ,n21[5]);
    not g2264(n388 ,n17[0]);
    not g2265(n387 ,n52[5]);
    not g2266(n386 ,n50[6]);
    not g2267(n385 ,n60[5]);
    not g2268(n384 ,n22[6]);
    not g2269(n383 ,n52[6]);
    not g2270(n382 ,n27[3]);
    not g2271(n381 ,n23[1]);
    not g2272(n380 ,n44[2]);
    not g2273(n379 ,n34[0]);
    not g2274(n378 ,n28[4]);
    not g2275(n377 ,n54[5]);
    not g2276(n376 ,n35[2]);
    not g2277(n375 ,n60[6]);
    not g2278(n374 ,n32[7]);
    not g2279(n373 ,n44[7]);
    not g2280(n372 ,n45[2]);
    not g2281(n371 ,n22[1]);
    not g2282(n370 ,n23[6]);
    not g2283(n369 ,n56[7]);
    not g2284(n368 ,n30[6]);
    not g2285(n367 ,n35[5]);
    not g2286(n366 ,n41[6]);
    not g2287(n365 ,n29[7]);
    not g2288(n364 ,n52[1]);
    not g2289(n363 ,n32[3]);
    not g2290(n362 ,n52[2]);
    not g2291(n361 ,n22[3]);
    not g2292(n360 ,n35[7]);
    not g2293(n359 ,n53[1]);
    not g2294(n358 ,n26[6]);
    not g2295(n357 ,n21[2]);
    not g2296(n356 ,n23[0]);
    not g2297(n355 ,n35[0]);
    not g2298(n354 ,n27[7]);
    not g2299(n353 ,n41[2]);
    not g2300(n352 ,n46[0]);
    not g2301(n351 ,n57[1]);
    not g2302(n350 ,n18[2]);
    not g2303(n349 ,n57[2]);
    not g2304(n348 ,n57[0]);
    not g2305(n347 ,n36[0]);
    not g2306(n346 ,n18[3]);
    not g2307(n345 ,n36[3]);
    not g2308(n344 ,n57[3]);
    not g2309(n343 ,n59[3]);
    not g2310(n342 ,n38[1]);
    not g2311(n341 ,n58[0]);
    not g2312(n340 ,n59[1]);
    not g2313(n339 ,n19[0]);
    not g2314(n338 ,n59[0]);
    not g2315(n337 ,n38[0]);
    not g2316(n336 ,n58[3]);
    not g2317(n335 ,n37[1]);
    not g2318(n334 ,n38[2]);
    not g2319(n333 ,n58[1]);
    not g2320(n332 ,n37[3]);
    not g2321(n331 ,n37[2]);
    not g2322(n330 ,n59[2]);
    not g2323(n329 ,n39[4]);
    not g2324(n328 ,n39[2]);
    not g2325(n327 ,n39[3]);
    not g2326(n326 ,n2310);
    not g2327(n325 ,n2305);
    not g2328(n324 ,n2324);
    not g2329(n323 ,n2320);
    not g2330(n322 ,n2309);
    not g2331(n321 ,n2300);
    not g2332(n320 ,n2303);
    not g2333(n319 ,n2327);
    not g2334(n318 ,n2325);
    not g2335(n317 ,n2326);
    not g2336(n316 ,n2331);
    not g2337(n315 ,n2329);
    not g2338(n314 ,n2307);
    not g2339(n313 ,n2306);
    not g2340(n312 ,n2323);
    not g2341(n311 ,n2328);
    not g2342(n310 ,n2301);
    not g2343(n309 ,n2313);
    not g2344(n308 ,n2304);
    not g2345(n307 ,n2314);
    not g2346(n306 ,n2321);
    not g2347(n305 ,n2317);
    not g2348(n304 ,n2302);
    not g2349(n303 ,n2318);
    not g2350(n302 ,n2308);
    not g2351(n301 ,n2315);
    not g2352(n300 ,n2322);
    not g2353(n299 ,n2330);
    not g2354(n298 ,n2319);
    not g2355(n297 ,n2311);
    not g2356(n296 ,n2312);
    not g2357(n295 ,n34[6]);
    not g2358(n294 ,n43[3]);
    not g2359(n293 ,n52[3]);
    not g2360(n292 ,n23[4]);
    not g2361(n291 ,n60[1]);
    not g2362(n290 ,n53[3]);
    not g2363(n289 ,n47[7]);
    not g2364(n288 ,n45[0]);
    not g2365(n287 ,n23[2]);
    not g2366(n286 ,n51[1]);
    not g2367(n285 ,n45[4]);
    not g2368(n284 ,n33[6]);
    not g2369(n283 ,n41[1]);
    not g2370(n282 ,n31[2]);
    not g2371(n281 ,n30[3]);
    not g2372(n280 ,n50[7]);
    not g2373(n279 ,n60[4]);
    not g2374(n278 ,n42[3]);
    not g2375(n277 ,n43[1]);
    not g2376(n276 ,n30[4]);
    not g2377(n275 ,n23[5]);
    not g2378(n274 ,n46[1]);
    not g2379(n273 ,n32[0]);
    not g2380(n272 ,n54[4]);
    not g2381(n271 ,n43[6]);
    not g2382(n270 ,n32[6]);
    not g2383(n269 ,n55[6]);
    not g2384(n268 ,n28[1]);
    not g2385(n267 ,n45[3]);
    not g2386(n266 ,n47[0]);
    not g2387(n265 ,n48[5]);
    not g2388(n264 ,n49[6]);
    not g2389(n263 ,n41[5]);
    not g2390(n262 ,n44[1]);
    not g2391(n261 ,n47[6]);
    not g2392(n260 ,n24[7]);
    not g2393(n259 ,n49[7]);
    not g2394(n258 ,n49[4]);
    not g2395(n257 ,n28[2]);
    not g2396(n256 ,n48[0]);
    not g2397(n255 ,n45[7]);
    not g2398(n254 ,n28[7]);
    not g2399(n253 ,n55[2]);
    not g2400(n252 ,n51[6]);
    not g2401(n251 ,n25[0]);
    not g2402(n250 ,n48[2]);
    not g2403(n249 ,n41[7]);
    not g2404(n248 ,n51[5]);
    not g2405(n247 ,n34[2]);
    not g2406(n246 ,n55[7]);
    not g2407(n245 ,n21[4]);
    not g2408(n244 ,n27[6]);
    not g2409(n243 ,n29[4]);
    not g2410(n242 ,n55[1]);
    not g2411(n241 ,n41[4]);
    not g2412(n240 ,n50[4]);
    not g2413(n239 ,n20[5]);
    not g2414(n238 ,n49[3]);
    not g2415(n237 ,n46[3]);
    not g2416(n236 ,n21[7]);
    not g2417(n235 ,n6[4]);
    not g2418(n234 ,n20[6]);
    not g2419(n233 ,n46[4]);
    not g2420(n232 ,n28[6]);
    not g2421(n231 ,n51[2]);
    not g2422(n230 ,n22[7]);
    not g2423(n229 ,n6[5]);
    not g2424(n228 ,n44[6]);
    not g2425(n227 ,n6[0]);
    not g2426(n226 ,n27[1]);
    not g2427(n225 ,n55[4]);
    not g2428(n224 ,n53[2]);
    not g2429(n223 ,n56[0]);
    not g2430(n222 ,n25[6]);
    not g2431(n221 ,n29[1]);
    not g2432(n220 ,n54[1]);
    not g2433(n219 ,n32[2]);
    not g2434(n218 ,n35[3]);
    not g2435(n217 ,n28[3]);
    not g2436(n216 ,n16);
    not g2437(n215 ,n42[5]);
    not g2438(n214 ,n34[1]);
    not g2439(n213 ,n45[5]);
    not g2440(n212 ,n50[0]);
    not g2441(n211 ,n8[1]);
    not g2442(n210 ,n53[4]);
    not g2443(n209 ,n31[5]);
    not g2444(n208 ,n20[2]);
    not g2445(n207 ,n53[6]);
    not g2446(n206 ,n43[4]);
    not g2447(n205 ,n33[7]);
    not g2448(n204 ,n26[7]);
    not g2449(n203 ,n33[5]);
    not g2450(n202 ,n24[5]);
    not g2451(n201 ,n50[3]);
    not g2452(n200 ,n60[0]);
    not g2453(n199 ,n49[1]);
    not g2454(n198 ,n17[3]);
    not g2455(n197 ,n29[0]);
    not g2456(n196 ,n6[2]);
    not g2457(n195 ,n24[0]);
    not g2458(n194 ,n30[1]);
    not g2459(n193 ,n32[4]);
    not g2460(n192 ,n6[7]);
    not g2461(n191 ,n33[4]);
    not g2462(n190 ,n42[0]);
    not g2463(n189 ,n6[1]);
    not g2464(n188 ,n2);
    not g2465(n187 ,n60[7]);
    not g2466(n186 ,n47[1]);
    not g2467(n185 ,n20[0]);
    not g2468(n184 ,n54[2]);
    not g2469(n183 ,n23[7]);
    not g2470(n182 ,n31[3]);
    not g2471(n181 ,n45[6]);
    not g2472(n180 ,n56[6]);
    not g2473(n179 ,n56[4]);
    not g2474(n178 ,n6[3]);
    not g2475(n177 ,n30[7]);
    not g2476(n176 ,n33[1]);
    not g2477(n175 ,n28[0]);
    not g2478(n174 ,n53[7]);
    not g2479(n173 ,n13);
    not g2480(n172 ,n19[1]);
    not g2481(n171 ,n36[2]);
    not g2482(n170 ,n18[1]);
    not g2483(n169 ,n36[1]);
    not g2484(n168 ,n18[0]);
    not g2485(n167 ,n37[0]);
    not g2486(n166 ,n38[3]);
    not g2487(n165 ,n15);
    not g2488(n164 ,n58[2]);
    not g2489(n163 ,n36[4]);
    not g2490(n162 ,n57[4]);
    not g2491(n161 ,n40[0]);
    not g2492(n160 ,n40[1]);
    not g2493(n159 ,n4[1]);
    not g2494(n158 ,n4[2]);
    not g2495(n157 ,n4[5]);
    not g2496(n156 ,n4[6]);
    not g2497(n155 ,n4[3]);
    not g2498(n154 ,n4[7]);
    not g2499(n153 ,n4[4]);
    not g2500(n152 ,n4[0]);
    not g2501(n151 ,n39[6]);
    not g2502(n150 ,n39[5]);
    not g2503(n149 ,n39[0]);
    not g2504(n148 ,n39[1]);
    not g2505(n147 ,n1);
    not g2506(n146 ,n1);
    not g2507(n145 ,n1);
    not g2508(n144 ,n1);
    not g2509(n143 ,n1);
    not g2510(n142 ,n1);
    not g2511(n141 ,n1);
    xor g2512(n2324 ,n57[4] ,n70);
    xor g2513(n2323 ,n57[3] ,n68);
    nor g2514(n70 ,n57[3] ,n69);
    xor g2515(n2322 ,n57[2] ,n66);
    not g2516(n69 ,n68);
    nor g2517(n68 ,n57[2] ,n67);
    xnor g2518(n2321 ,n57[1] ,n57[0]);
    not g2519(n67 ,n66);
    nor g2520(n66 ,n57[1] ,n57[0]);
    xor g2521(n2312 ,n36[4] ,n65);
    xor g2522(n2327 ,n36[3] ,n63);
    nor g2523(n65 ,n36[3] ,n64);
    xor g2524(n2326 ,n36[2] ,n61);
    not g2525(n64 ,n63);
    nor g2526(n63 ,n36[2] ,n62);
    xnor g2527(n2325 ,n36[1] ,n36[0]);
    not g2528(n62 ,n61);
    nor g2529(n61 ,n36[1] ,n36[0]);
    or g2530(n2333 ,n72 ,n73);
    or g2531(n73 ,n57[3] ,n71);
    or g2532(n72 ,n57[2] ,n57[0]);
    or g2533(n71 ,n57[4] ,n57[1]);
    or g2534(n2332 ,n75 ,n76);
    or g2535(n76 ,n36[3] ,n74);
    or g2536(n75 ,n36[2] ,n36[0]);
    or g2537(n74 ,n36[4] ,n36[1]);
    xor g2538(n2320 ,n57[4] ,n100);
    nor g2539(n2319 ,n99 ,n100);
    nor g2540(n100 ,n90 ,n98);
    nor g2541(n99 ,n57[3] ,n97);
    nor g2542(n2318 ,n96 ,n97);
    not g2543(n98 ,n97);
    nor g2544(n97 ,n92 ,n95);
    nor g2545(n96 ,n57[2] ,n94);
    nor g2546(n2317 ,n94 ,n93);
    not g2547(n95 ,n94);
    nor g2548(n94 ,n89 ,n91);
    nor g2549(n93 ,n57[1] ,n57[0]);
    not g2550(n92 ,n57[2]);
    not g2551(n91 ,n57[0]);
    not g2552(n90 ,n57[3]);
    not g2553(n89 ,n57[1]);
    nor g2554(n2314 ,n87 ,n88);
    nor g2555(n88 ,n78 ,n86);
    nor g2556(n87 ,n36[3] ,n85);
    nor g2557(n2313 ,n84 ,n85);
    not g2558(n86 ,n85);
    nor g2559(n85 ,n80 ,n83);
    nor g2560(n84 ,n36[2] ,n82);
    nor g2561(n2328 ,n82 ,n81);
    not g2562(n83 ,n82);
    nor g2563(n82 ,n77 ,n79);
    nor g2564(n81 ,n36[1] ,n36[0]);
    not g2565(n80 ,n36[2]);
    not g2566(n79 ,n36[0]);
    not g2567(n78 ,n36[3]);
    not g2568(n77 ,n36[1]);
    xor g2569(n2302 ,n59[3] ,n108);
    nor g2570(n2301 ,n107 ,n108);
    nor g2571(n108 ,n103 ,n106);
    nor g2572(n107 ,n59[2] ,n105);
    nor g2573(n2300 ,n105 ,n104);
    not g2574(n106 ,n105);
    nor g2575(n105 ,n101 ,n102);
    nor g2576(n104 ,n59[1] ,n59[0]);
    not g2577(n103 ,n59[2]);
    not g2578(n102 ,n59[0]);
    not g2579(n101 ,n59[1]);
    xor g2580(n2305 ,n37[3] ,n116);
    nor g2581(n2304 ,n115 ,n116);
    nor g2582(n116 ,n111 ,n114);
    nor g2583(n115 ,n37[2] ,n113);
    nor g2584(n2303 ,n113 ,n112);
    not g2585(n114 ,n113);
    nor g2586(n113 ,n109 ,n110);
    nor g2587(n112 ,n37[1] ,n37[0]);
    not g2588(n111 ,n37[2]);
    not g2589(n110 ,n37[0]);
    not g2590(n109 ,n37[1]);
    xor g2591(n2308 ,n58[3] ,n124);
    nor g2592(n2307 ,n123 ,n124);
    nor g2593(n124 ,n119 ,n122);
    nor g2594(n123 ,n58[2] ,n121);
    nor g2595(n2306 ,n121 ,n120);
    not g2596(n122 ,n121);
    nor g2597(n121 ,n117 ,n118);
    nor g2598(n120 ,n58[1] ,n58[0]);
    not g2599(n119 ,n58[2]);
    not g2600(n118 ,n58[0]);
    not g2601(n117 ,n58[1]);
    xor g2602(n2316 ,n19[1] ,n19[0]);
    xor g2603(n2311 ,n38[3] ,n132);
    nor g2604(n2310 ,n131 ,n132);
    nor g2605(n132 ,n127 ,n130);
    nor g2606(n131 ,n38[2] ,n129);
    nor g2607(n2309 ,n129 ,n128);
    not g2608(n130 ,n129);
    nor g2609(n129 ,n125 ,n126);
    nor g2610(n128 ,n38[1] ,n38[0]);
    not g2611(n127 ,n38[2]);
    not g2612(n126 ,n38[0]);
    not g2613(n125 ,n38[1]);
    xor g2614(n2331 ,n18[3] ,n140);
    nor g2615(n2330 ,n139 ,n140);
    nor g2616(n140 ,n135 ,n138);
    nor g2617(n139 ,n18[2] ,n137);
    nor g2618(n2329 ,n137 ,n136);
    not g2619(n138 ,n137);
    nor g2620(n137 ,n133 ,n134);
    nor g2621(n136 ,n18[1] ,n18[0]);
    not g2622(n135 ,n18[2]);
    not g2623(n134 ,n18[0]);
    not g2624(n133 ,n18[1]);
    buf g2625(n580 ,n557);
    buf g2626(n2315 ,n88);
    not g2627(n1004 ,n554);
endmodule
