module top(n0, n1, n2, n6, n3, n7, n5, n12, n4, n8, n9, n10, n11, n13, n14, n15, n16);
    input n0, n1, n2, n3, n4;
    input [7:0] n5;
    output n6, n7, n8, n9, n10, n11;
    output [7:0] n12, n13, n14, n15;
    output [15:0] n16;
    wire n0, n1, n2, n3, n4;
    wire [7:0] n5;
    wire n6, n7, n8, n9, n10, n11;
    wire [7:0] n12, n13, n14, n15;
    wire [15:0] n16;
    wire [2:0] n17;
    wire [2:0] n18;
    wire [4:0] n19;
    wire [15:0] n20;
    wire [7:0] n21;
    wire [7:0] n22;
    wire [7:0] n23;
    wire [7:0] n24;
    wire [7:0] n25;
    wire [7:0] n26;
    wire [7:0] n27;
    wire [7:0] n28;
    wire [7:0] n29;
    wire [7:0] n30;
    wire [7:0] n31;
    wire [7:0] n32;
    wire [7:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [7:0] n36;
    wire [3:0] n37;
    wire [3:0] n38;
    wire [7:0] n39;
    wire [15:0] n40;
    wire [2:0] n41;
    wire [7:0] n42;
    wire [7:0] n43;
    wire [7:0] n44;
    wire [7:0] n45;
    wire [7:0] n46;
    wire [7:0] n47;
    wire [7:0] n48;
    wire [7:0] n49;
    wire [7:0] n50;
    wire [7:0] n51;
    wire [7:0] n52;
    wire [7:0] n53;
    wire [7:0] n54;
    wire [7:0] n55;
    wire [7:0] n56;
    wire [7:0] n57;
    wire [4:0] n58;
    wire [3:0] n59;
    wire [3:0] n60;
    wire [7:0] n61;
    wire [2:0] n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848, n849, n850, n851, n852, n853, n854;
    wire n855, n856, n857, n858, n859, n860, n861, n862;
    wire n863, n864, n865, n866, n867, n868, n869, n870;
    wire n871, n872, n873, n874, n875, n876, n877, n878;
    wire n879, n880, n881, n882, n883, n884, n885, n886;
    wire n887, n888, n889, n890, n891, n892, n893, n894;
    wire n895, n896, n897, n898, n899, n900, n901, n902;
    wire n903, n904, n905, n906, n907, n908, n909, n910;
    wire n911, n912, n913, n914, n915, n916, n917, n918;
    wire n919, n920, n921, n922, n923, n924, n925, n926;
    wire n927, n928, n929, n930, n931, n932, n933, n934;
    wire n935, n936, n937, n938, n939, n940, n941, n942;
    wire n943, n944, n945, n946, n947, n948, n949, n950;
    wire n951, n952, n953, n954, n955, n956, n957, n958;
    wire n959, n960, n961, n962, n963, n964, n965, n966;
    wire n967, n968, n969, n970, n971, n972, n973, n974;
    wire n975, n976, n977, n978, n979, n980, n981, n982;
    wire n983, n984, n985, n986, n987, n988, n989, n990;
    wire n991, n992, n993, n994, n995, n996, n997, n998;
    wire n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
    wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
    wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
    wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
    wire n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
    wire n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
    wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
    wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
    wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
    wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
    wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
    wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
    wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
    wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
    wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
    wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
    wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
    wire n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142;
    wire n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
    wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158;
    wire n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166;
    wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
    wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
    wire n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190;
    wire n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198;
    wire n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206;
    wire n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
    wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
    wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
    wire n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238;
    wire n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246;
    wire n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254;
    wire n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;
    wire n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;
    wire n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;
    wire n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;
    wire n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;
    wire n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;
    wire n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;
    wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
    wire n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;
    wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
    wire n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;
    wire n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;
    wire n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;
    wire n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;
    wire n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;
    wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
    wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
    wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
    wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
    wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
    wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
    wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
    wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
    wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
    wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
    wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
    wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
    wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
    wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
    wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
    wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
    wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
    wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
    wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
    wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
    wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
    wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
    wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
    wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
    wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
    wire n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582;
    wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
    wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
    wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
    wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
    wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
    wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
    wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
    wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
    wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
    wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
    wire n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
    wire n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678;
    wire n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686;
    wire n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694;
    wire n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702;
    wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
    wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
    wire n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726;
    wire n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734;
    wire n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742;
    wire n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750;
    wire n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758;
    wire n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766;
    wire n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774;
    wire n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782;
    wire n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790;
    wire n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798;
    wire n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806;
    wire n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814;
    wire n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822;
    wire n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;
    wire n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838;
    wire n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846;
    wire n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854;
    wire n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862;
    wire n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870;
    wire n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878;
    wire n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886;
    wire n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894;
    wire n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902;
    wire n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910;
    wire n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918;
    wire n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926;
    wire n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934;
    wire n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942;
    wire n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950;
    wire n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958;
    wire n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966;
    wire n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974;
    wire n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982;
    wire n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990;
    wire n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998;
    wire n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006;
    wire n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014;
    wire n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022;
    wire n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030;
    wire n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038;
    wire n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046;
    wire n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054;
    wire n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062;
    wire n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070;
    wire n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078;
    wire n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086;
    wire n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094;
    wire n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102;
    wire n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110;
    wire n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118;
    wire n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126;
    wire n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134;
    wire n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142;
    wire n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150;
    wire n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158;
    wire n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166;
    wire n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174;
    wire n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182;
    wire n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190;
    wire n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198;
    wire n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206;
    wire n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214;
    wire n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222;
    wire n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230;
    wire n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238;
    wire n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246;
    wire n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254;
    wire n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262;
    wire n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270;
    wire n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278;
    wire n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286;
    wire n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294;
    wire n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302;
    wire n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310;
    wire n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318;
    wire n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326;
    wire n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334;
    wire n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342;
    wire n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350;
    wire n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358;
    wire n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366;
    wire n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374;
    wire n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382;
    wire n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390;
    wire n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398;
    wire n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406;
    wire n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414;
    wire n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422;
    wire n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430;
    wire n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438;
    wire n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446;
    wire n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454;
    wire n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462;
    wire n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470;
    wire n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478;
    wire n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486;
    wire n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494;
    wire n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502;
    wire n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510;
    wire n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518;
    wire n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526;
    wire n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534;
    wire n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542;
    wire n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550;
    wire n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558;
    wire n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566;
    wire n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574;
    wire n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582;
    wire n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590;
    wire n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598;
    wire n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606;
    wire n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614;
    wire n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622;
    wire n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630;
    wire n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638;
    wire n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646;
    wire n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654;
    wire n2655;
    buf g0(n16[11], 1'b0);
    buf g1(n16[12], 1'b0);
    buf g2(n16[13], 1'b0);
    buf g3(n16[14], 1'b0);
    buf g4(n16[15], 1'b0);
    buf g5(n15[0], 1'b0);
    buf g6(n15[1], 1'b0);
    buf g7(n15[2], 1'b0);
    buf g8(n15[3], n13[1]);
    buf g9(n15[4], n13[2]);
    buf g10(n15[5], n13[5]);
    buf g11(n14[0], 1'b0);
    buf g12(n14[2], 1'b0);
    buf g13(n14[3], 1'b0);
    buf g14(n14[4], 1'b0);
    buf g15(n14[5], 1'b0);
    buf g16(n14[6], 1'b0);
    buf g17(n14[7], 1'b0);
    buf g18(n13[0], 1'b0);
    not g19(n2597 ,n2647);
    not g20(n2596 ,n2621);
    not g21(n2595 ,n17[2]);
    or g22(n2618 ,n2592 ,n2594);
    or g23(n2594 ,n2591 ,n2593);
    or g24(n2593 ,n2589 ,n2646);
    or g25(n2646 ,n18[0] ,n2590);
    or g26(n2592 ,n2595 ,n17[1]);
    or g27(n2591 ,n19[4] ,n17[0]);
    or g28(n2590 ,n18[2] ,n18[1]);
    not g29(n2589 ,n2654);
    dff g30(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n743), .Q(n16[0]));
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n731), .Q(n16[1]));
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n740), .Q(n16[2]));
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n737), .Q(n16[3]));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n742), .Q(n16[4]));
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n732), .Q(n16[5]));
    dff g36(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n738), .Q(n16[6]));
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n735), .Q(n16[7]));
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n733), .Q(n16[8]));
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n739), .Q(n16[9]));
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n734), .Q(n16[10]));
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n700), .Q(n7));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1780), .Q(n14[1]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n759), .Q(n13[1]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n898), .Q(n13[2]));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n871), .Q(n13[5]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n741), .Q(n15[6]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n730), .Q(n15[7]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2341), .Q(n20[0]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2338), .Q(n20[1]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2355), .Q(n20[2]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2345), .Q(n20[3]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2340), .Q(n20[4]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2466), .Q(n20[5]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2458), .Q(n20[6]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2464), .Q(n20[7]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2460), .Q(n20[8]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2451), .Q(n20[9]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2448), .Q(n20[10]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2445), .Q(n20[11]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2437), .Q(n20[12]));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2028), .Q(n18[0]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2021), .Q(n18[1]));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2010), .Q(n18[2]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1814), .Q(n11));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2535), .Q(n12[0]));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2537), .Q(n12[1]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2536), .Q(n12[2]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2534), .Q(n12[3]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2546), .Q(n12[4]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2545), .Q(n12[5]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2539), .Q(n12[6]));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2538), .Q(n12[7]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1819), .Q(n9));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2399), .Q(n21[0]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2397), .Q(n21[1]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2398), .Q(n21[2]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2396), .Q(n21[3]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2395), .Q(n21[4]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2394), .Q(n21[5]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2393), .Q(n21[6]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2392), .Q(n21[7]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2391), .Q(n22[0]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2390), .Q(n22[1]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2389), .Q(n22[2]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2388), .Q(n22[3]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2387), .Q(n22[4]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2386), .Q(n22[5]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2384), .Q(n22[6]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2385), .Q(n22[7]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2383), .Q(n23[0]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2382), .Q(n23[1]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2381), .Q(n23[2]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2380), .Q(n23[3]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2379), .Q(n23[4]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2378), .Q(n23[5]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2377), .Q(n23[6]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2376), .Q(n23[7]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2375), .Q(n24[0]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2374), .Q(n24[1]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2373), .Q(n24[2]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2372), .Q(n24[3]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2371), .Q(n24[4]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2370), .Q(n24[5]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2369), .Q(n24[6]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2368), .Q(n24[7]));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2367), .Q(n25[0]));
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2366), .Q(n25[1]));
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2365), .Q(n25[2]));
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2364), .Q(n25[3]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2363), .Q(n25[4]));
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2362), .Q(n25[5]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2361), .Q(n25[6]));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2360), .Q(n25[7]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2359), .Q(n26[0]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2358), .Q(n26[1]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2357), .Q(n26[2]));
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2356), .Q(n26[3]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2354), .Q(n26[4]));
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2353), .Q(n26[5]));
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2352), .Q(n26[6]));
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2351), .Q(n26[7]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2350), .Q(n27[0]));
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2349), .Q(n27[1]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2348), .Q(n27[2]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2347), .Q(n27[3]));
    dff g126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2346), .Q(n27[4]));
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2344), .Q(n27[5]));
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2343), .Q(n27[6]));
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2342), .Q(n27[7]));
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2339), .Q(n28[0]));
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2337), .Q(n28[1]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2336), .Q(n28[2]));
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2474), .Q(n28[3]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2473), .Q(n28[4]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2514), .Q(n28[5]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2471), .Q(n28[6]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2470), .Q(n28[7]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2469), .Q(n29[0]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2468), .Q(n29[1]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2467), .Q(n29[2]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2465), .Q(n29[3]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2463), .Q(n29[4]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2462), .Q(n29[5]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2461), .Q(n29[6]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2459), .Q(n29[7]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2457), .Q(n30[0]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2456), .Q(n30[1]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2455), .Q(n30[2]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2454), .Q(n30[3]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2453), .Q(n30[4]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2452), .Q(n30[5]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2450), .Q(n30[6]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2449), .Q(n30[7]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2447), .Q(n31[0]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2446), .Q(n31[1]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2444), .Q(n31[2]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2443), .Q(n31[3]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2442), .Q(n31[4]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2440), .Q(n31[5]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2436), .Q(n31[6]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2435), .Q(n31[7]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2434), .Q(n32[0]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2433), .Q(n32[1]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2432), .Q(n32[2]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2431), .Q(n32[3]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2430), .Q(n32[4]));
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2510), .Q(n32[5]));
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2511), .Q(n32[6]));
    dff g169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2512), .Q(n32[7]));
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2513), .Q(n33[0]));
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2472), .Q(n33[1]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2429), .Q(n33[2]));
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2428), .Q(n33[3]));
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2427), .Q(n33[4]));
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2426), .Q(n33[5]));
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2425), .Q(n33[6]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2424), .Q(n33[7]));
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2423), .Q(n34[0]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2422), .Q(n34[1]));
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2421), .Q(n34[2]));
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2420), .Q(n34[3]));
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2419), .Q(n34[4]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2418), .Q(n34[5]));
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2417), .Q(n34[6]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2416), .Q(n34[7]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2415), .Q(n35[0]));
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2413), .Q(n35[1]));
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2414), .Q(n35[2]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2412), .Q(n35[3]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2411), .Q(n35[4]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2410), .Q(n35[5]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2409), .Q(n35[6]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2408), .Q(n35[7]));
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2407), .Q(n36[0]));
    dff g195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2406), .Q(n36[1]));
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2405), .Q(n36[2]));
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2404), .Q(n36[3]));
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2403), .Q(n36[4]));
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2402), .Q(n36[5]));
    dff g200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2401), .Q(n36[6]));
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2400), .Q(n36[7]));
    dff g202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1813), .Q(n19[0]));
    dff g203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1815), .Q(n19[1]));
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1816), .Q(n19[2]));
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1817), .Q(n19[3]));
    dff g206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1818), .Q(n19[4]));
    dff g207(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n815), .Q(n37[0]));
    dff g208(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1618), .Q(n37[1]));
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1617), .Q(n37[2]));
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1616), .Q(n37[3]));
    dff g211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1774), .Q(n38[0]));
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2515), .Q(n38[1]));
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2517), .Q(n38[2]));
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2516), .Q(n38[3]));
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n936), .Q(n39[0]));
    dff g216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n937), .Q(n39[1]));
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n935), .Q(n39[2]));
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n938), .Q(n39[3]));
    dff g219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n941), .Q(n39[4]));
    dff g220(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n939), .Q(n39[5]));
    dff g221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n942), .Q(n39[6]));
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n940), .Q(n39[7]));
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2051), .Q(n17[0]));
    dff g224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2050), .Q(n17[1]));
    dff g225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2049), .Q(n17[2]));
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n913), .Q(n13[3]));
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n872), .Q(n13[4]));
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n744), .Q(n13[6]));
    dff g229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n736), .Q(n13[7]));
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1659), .Q(n40[0]));
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1658), .Q(n40[1]));
    dff g232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1657), .Q(n40[2]));
    dff g233(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1656), .Q(n40[3]));
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1655), .Q(n40[4]));
    dff g235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1654), .Q(n40[5]));
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1653), .Q(n40[6]));
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1652), .Q(n40[7]));
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1651), .Q(n40[8]));
    dff g239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1650), .Q(n40[9]));
    dff g240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1649), .Q(n40[10]));
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1776), .Q(n41[0]));
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1778), .Q(n41[1]));
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1779), .Q(n41[2]));
    dff g244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1765), .Q(n10));
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1766), .Q(n8));
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1611), .Q(n42[0]));
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1610), .Q(n42[1]));
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1609), .Q(n42[2]));
    dff g249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1608), .Q(n42[3]));
    dff g250(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1607), .Q(n42[4]));
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1606), .Q(n42[5]));
    dff g252(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1605), .Q(n42[6]));
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1604), .Q(n42[7]));
    dff g254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1603), .Q(n43[0]));
    dff g255(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1602), .Q(n43[1]));
    dff g256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1601), .Q(n43[2]));
    dff g257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1600), .Q(n43[3]));
    dff g258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1599), .Q(n43[4]));
    dff g259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1598), .Q(n43[5]));
    dff g260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1597), .Q(n43[6]));
    dff g261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1596), .Q(n43[7]));
    dff g262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1595), .Q(n44[0]));
    dff g263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1594), .Q(n44[1]));
    dff g264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1593), .Q(n44[2]));
    dff g265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1592), .Q(n44[3]));
    dff g266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1591), .Q(n44[4]));
    dff g267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1590), .Q(n44[5]));
    dff g268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1589), .Q(n44[6]));
    dff g269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1588), .Q(n44[7]));
    dff g270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1587), .Q(n45[0]));
    dff g271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1586), .Q(n45[1]));
    dff g272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1585), .Q(n45[2]));
    dff g273(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1584), .Q(n45[3]));
    dff g274(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1583), .Q(n45[4]));
    dff g275(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1621), .Q(n45[5]));
    dff g276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1581), .Q(n45[6]));
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1580), .Q(n45[7]));
    dff g278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1579), .Q(n46[0]));
    dff g279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1578), .Q(n46[1]));
    dff g280(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1577), .Q(n46[2]));
    dff g281(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1576), .Q(n46[3]));
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1575), .Q(n46[4]));
    dff g283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1574), .Q(n46[5]));
    dff g284(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1573), .Q(n46[6]));
    dff g285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1572), .Q(n46[7]));
    dff g286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1571), .Q(n47[0]));
    dff g287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1569), .Q(n47[1]));
    dff g288(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1568), .Q(n47[2]));
    dff g289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1567), .Q(n47[3]));
    dff g290(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1566), .Q(n47[4]));
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1565), .Q(n47[5]));
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1564), .Q(n47[6]));
    dff g293(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1563), .Q(n47[7]));
    dff g294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1562), .Q(n48[0]));
    dff g295(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1561), .Q(n48[1]));
    dff g296(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1560), .Q(n48[2]));
    dff g297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1559), .Q(n48[3]));
    dff g298(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1558), .Q(n48[4]));
    dff g299(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1622), .Q(n48[5]));
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1556), .Q(n48[6]));
    dff g301(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1555), .Q(n48[7]));
    dff g302(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1554), .Q(n49[0]));
    dff g303(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1553), .Q(n49[1]));
    dff g304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1552), .Q(n49[2]));
    dff g305(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1551), .Q(n49[3]));
    dff g306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1550), .Q(n49[4]));
    dff g307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1549), .Q(n49[5]));
    dff g308(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1548), .Q(n49[6]));
    dff g309(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1547), .Q(n49[7]));
    dff g310(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1546), .Q(n50[0]));
    dff g311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1545), .Q(n50[1]));
    dff g312(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1544), .Q(n50[2]));
    dff g313(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1543), .Q(n50[3]));
    dff g314(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1542), .Q(n50[4]));
    dff g315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1541), .Q(n50[5]));
    dff g316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1540), .Q(n50[6]));
    dff g317(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1539), .Q(n50[7]));
    dff g318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1538), .Q(n51[0]));
    dff g319(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1537), .Q(n51[1]));
    dff g320(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1536), .Q(n51[2]));
    dff g321(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1535), .Q(n51[3]));
    dff g322(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1534), .Q(n51[4]));
    dff g323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1533), .Q(n51[5]));
    dff g324(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1532), .Q(n51[6]));
    dff g325(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1531), .Q(n51[7]));
    dff g326(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1582), .Q(n52[0]));
    dff g327(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1529), .Q(n52[1]));
    dff g328(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1528), .Q(n52[2]));
    dff g329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1620), .Q(n52[3]));
    dff g330(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1527), .Q(n52[4]));
    dff g331(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1526), .Q(n52[5]));
    dff g332(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1525), .Q(n52[6]));
    dff g333(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1524), .Q(n52[7]));
    dff g334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1522), .Q(n53[0]));
    dff g335(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1521), .Q(n53[1]));
    dff g336(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1520), .Q(n53[2]));
    dff g337(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1519), .Q(n53[3]));
    dff g338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1518), .Q(n53[4]));
    dff g339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1517), .Q(n53[5]));
    dff g340(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1614), .Q(n53[6]));
    dff g341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1648), .Q(n53[7]));
    dff g342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1647), .Q(n54[0]));
    dff g343(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1646), .Q(n54[1]));
    dff g344(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1645), .Q(n54[2]));
    dff g345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1644), .Q(n54[3]));
    dff g346(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1643), .Q(n54[4]));
    dff g347(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1642), .Q(n54[5]));
    dff g348(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1641), .Q(n54[6]));
    dff g349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1640), .Q(n54[7]));
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1625), .Q(n55[0]));
    dff g351(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1639), .Q(n55[1]));
    dff g352(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1638), .Q(n55[2]));
    dff g353(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1637), .Q(n55[3]));
    dff g354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1636), .Q(n55[4]));
    dff g355(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1635), .Q(n55[5]));
    dff g356(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1619), .Q(n55[6]));
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1634), .Q(n55[7]));
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1633), .Q(n56[0]));
    dff g359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1632), .Q(n56[1]));
    dff g360(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1631), .Q(n56[2]));
    dff g361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1630), .Q(n56[3]));
    dff g362(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1629), .Q(n56[4]));
    dff g363(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1623), .Q(n56[5]));
    dff g364(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1628), .Q(n56[6]));
    dff g365(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1661), .Q(n56[7]));
    dff g366(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1662), .Q(n57[0]));
    dff g367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1664), .Q(n57[1]));
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1667), .Q(n57[2]));
    dff g369(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1668), .Q(n57[3]));
    dff g370(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1673), .Q(n57[4]));
    dff g371(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1699), .Q(n57[5]));
    dff g372(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1615), .Q(n57[6]));
    dff g373(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1700), .Q(n57[7]));
    dff g374(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1523), .Q(n58[0]));
    dff g375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1764), .Q(n58[1]));
    dff g376(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1755), .Q(n58[2]));
    dff g377(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1756), .Q(n58[3]));
    dff g378(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1757), .Q(n58[4]));
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1660), .Q(n59[0]));
    dff g380(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2441), .Q(n59[1]));
    dff g381(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2439), .Q(n59[2]));
    dff g382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2438), .Q(n59[3]));
    dff g383(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n880), .Q(n60[0]));
    dff g384(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1768), .Q(n60[1]));
    dff g385(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1770), .Q(n60[2]));
    dff g386(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1769), .Q(n60[3]));
    dff g387(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1345), .Q(n6));
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2585), .Q(n61[0]));
    dff g389(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2588), .Q(n61[1]));
    dff g390(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2587), .Q(n61[2]));
    dff g391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2586), .Q(n61[3]));
    dff g392(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2583), .Q(n61[4]));
    dff g393(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2584), .Q(n61[5]));
    dff g394(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2582), .Q(n61[6]));
    dff g395(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2574), .Q(n61[7]));
    dff g396(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2054), .Q(n62[0]));
    dff g397(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2053), .Q(n62[1]));
    dff g398(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2052), .Q(n62[2]));
    or g399(n2588 ,n1830 ,n2580);
    or g400(n2587 ,n1828 ,n2581);
    or g401(n2586 ,n1829 ,n2578);
    or g402(n2585 ,n1877 ,n2579);
    or g403(n2584 ,n1832 ,n2576);
    or g404(n2583 ,n1826 ,n2575);
    or g405(n2582 ,n1833 ,n2577);
    or g406(n2581 ,n969 ,n2573);
    or g407(n2580 ,n1115 ,n2572);
    or g408(n2579 ,n1105 ,n2571);
    or g409(n2578 ,n1091 ,n2570);
    or g410(n2577 ,n1078 ,n2569);
    or g411(n2576 ,n1098 ,n2568);
    or g412(n2575 ,n1133 ,n2567);
    or g413(n2574 ,n1868 ,n2566);
    or g414(n2573 ,n1853 ,n2565);
    or g415(n2572 ,n1941 ,n2564);
    or g416(n2571 ,n1956 ,n2563);
    or g417(n2570 ,n1839 ,n2562);
    or g418(n2569 ,n1971 ,n2561);
    or g419(n2568 ,n1930 ,n2560);
    or g420(n2567 ,n1914 ,n2559);
    or g421(n2566 ,n1827 ,n2558);
    or g422(n2565 ,n2498 ,n2555);
    or g423(n2564 ,n2501 ,n2556);
    or g424(n2563 ,n2504 ,n2553);
    or g425(n2562 ,n2494 ,n2554);
    or g426(n2561 ,n2485 ,n2551);
    or g427(n2560 ,n2488 ,n2552);
    or g428(n2559 ,n2491 ,n2557);
    or g429(n2558 ,n2482 ,n2550);
    or g430(n2557 ,n2012 ,n2543);
    or g431(n2556 ,n2033 ,n2547);
    or g432(n2555 ,n2026 ,n2548);
    or g433(n2554 ,n2020 ,n2549);
    or g434(n2553 ,n2041 ,n2544);
    or g435(n2552 ,n2005 ,n2542);
    or g436(n2551 ,n2000 ,n2541);
    or g437(n2550 ,n1995 ,n2540);
    or g438(n2549 ,n1852 ,n2530);
    or g439(n2548 ,n1926 ,n2531);
    or g440(n2547 ,n1921 ,n2532);
    or g441(n2546 ,n979 ,n2525);
    or g442(n2545 ,n1129 ,n2533);
    or g443(n2544 ,n1963 ,n2524);
    or g444(n2543 ,n1943 ,n2529);
    or g445(n2542 ,n1983 ,n2528);
    or g446(n2541 ,n1872 ,n2527);
    or g447(n2540 ,n1874 ,n2526);
    or g448(n2539 ,n1112 ,n2522);
    or g449(n2538 ,n1062 ,n2521);
    or g450(n2537 ,n984 ,n2520);
    or g451(n2536 ,n1125 ,n2519);
    or g452(n2535 ,n1101 ,n2523);
    or g453(n2534 ,n1132 ,n2518);
    or g454(n2533 ,n965 ,n2495);
    or g455(n2532 ,n2500 ,n2499);
    or g456(n2531 ,n2497 ,n2496);
    or g457(n2530 ,n2493 ,n2492);
    or g458(n2529 ,n2490 ,n2489);
    or g459(n2528 ,n2487 ,n2486);
    or g460(n2527 ,n2484 ,n2483);
    or g461(n2526 ,n2481 ,n2480);
    or g462(n2525 ,n959 ,n2505);
    or g463(n2524 ,n2503 ,n2502);
    or g464(n2523 ,n962 ,n2478);
    or g465(n2522 ,n963 ,n2479);
    or g466(n2521 ,n961 ,n2477);
    or g467(n2520 ,n960 ,n2476);
    or g468(n2519 ,n964 ,n2475);
    or g469(n2518 ,n966 ,n2506);
    or g470(n2517 ,n1696 ,n2509);
    or g471(n2516 ,n1695 ,n2507);
    or g472(n2515 ,n1697 ,n2508);
    or g473(n2514 ,n2311 ,n2055);
    or g474(n2513 ,n2275 ,n2173);
    or g475(n2512 ,n2276 ,n2135);
    or g476(n2511 ,n2277 ,n2136);
    or g477(n2510 ,n2278 ,n2137);
    nor g478(n2509 ,n465 ,n2166);
    nor g479(n2508 ,n461 ,n2166);
    nor g480(n2507 ,n478 ,n2166);
    or g481(n2506 ,n1694 ,n2185);
    or g482(n2505 ,n1678 ,n2184);
    or g483(n2504 ,n2043 ,n2042);
    or g484(n2503 ,n2039 ,n2038);
    or g485(n2502 ,n2037 ,n2036);
    or g486(n2501 ,n2035 ,n2034);
    or g487(n2500 ,n2032 ,n2031);
    or g488(n2499 ,n1992 ,n2030);
    or g489(n2498 ,n1990 ,n2027);
    or g490(n2497 ,n2025 ,n2024);
    or g491(n2496 ,n2023 ,n2165);
    or g492(n2495 ,n1674 ,n2183);
    or g493(n2494 ,n2022 ,n1991);
    or g494(n2493 ,n2019 ,n2018);
    or g495(n2492 ,n2017 ,n2016);
    or g496(n2491 ,n2014 ,n2013);
    or g497(n2490 ,n2011 ,n2009);
    or g498(n2489 ,n2007 ,n2008);
    or g499(n2488 ,n2029 ,n2006);
    or g500(n2487 ,n2004 ,n2044);
    or g501(n2486 ,n2045 ,n2046);
    or g502(n2485 ,n2002 ,n2001);
    or g503(n2484 ,n2047 ,n1999);
    or g504(n2483 ,n1998 ,n1997);
    or g505(n2482 ,n2015 ,n1996);
    or g506(n2481 ,n2040 ,n2003);
    or g507(n2480 ,n1994 ,n1993);
    or g508(n2479 ,n1689 ,n2182);
    or g509(n2478 ,n1688 ,n2181);
    or g510(n2477 ,n1685 ,n2180);
    or g511(n2476 ,n1679 ,n2179);
    or g512(n2475 ,n1727 ,n2178);
    or g513(n2474 ,n2313 ,n2333);
    or g514(n2473 ,n2312 ,n2334);
    or g515(n2472 ,n2274 ,n2134);
    or g516(n2471 ,n2310 ,n2164);
    or g517(n2470 ,n2309 ,n2163);
    or g518(n2469 ,n2308 ,n2177);
    or g519(n2468 ,n2307 ,n2162);
    or g520(n2467 ,n2306 ,n2161);
    or g521(n2466 ,n1490 ,n2325);
    or g522(n2465 ,n2305 ,n2160);
    or g523(n2464 ,n1484 ,n2323);
    or g524(n2463 ,n2304 ,n2159);
    or g525(n2462 ,n2303 ,n2158);
    or g526(n2461 ,n2302 ,n2157);
    or g527(n2460 ,n1488 ,n2322);
    or g528(n2459 ,n2301 ,n2156);
    or g529(n2458 ,n1489 ,n2324);
    or g530(n2457 ,n2300 ,n2176);
    or g531(n2456 ,n2299 ,n2155);
    or g532(n2455 ,n2298 ,n2154);
    or g533(n2454 ,n2297 ,n2153);
    or g534(n2453 ,n2296 ,n2152);
    or g535(n2452 ,n2295 ,n2151);
    or g536(n2451 ,n1487 ,n2321);
    or g537(n2450 ,n2294 ,n2150);
    or g538(n2449 ,n2293 ,n2149);
    or g539(n2448 ,n1480 ,n2320);
    or g540(n2447 ,n2292 ,n2175);
    or g541(n2446 ,n2291 ,n2148);
    or g542(n2445 ,n1483 ,n2319);
    or g543(n2444 ,n2290 ,n2147);
    or g544(n2443 ,n2289 ,n2146);
    or g545(n2442 ,n2288 ,n2145);
    or g546(n2441 ,n1349 ,n2328);
    or g547(n2440 ,n2287 ,n2144);
    or g548(n2439 ,n1348 ,n2327);
    or g549(n2438 ,n1500 ,n2326);
    or g550(n2437 ,n1486 ,n2318);
    or g551(n2436 ,n2286 ,n2143);
    or g552(n2435 ,n2285 ,n2142);
    or g553(n2434 ,n2284 ,n2174);
    or g554(n2433 ,n2283 ,n2141);
    or g555(n2432 ,n2282 ,n2140);
    or g556(n2431 ,n2281 ,n2139);
    or g557(n2430 ,n2279 ,n2138);
    or g558(n2429 ,n2273 ,n2133);
    or g559(n2428 ,n2272 ,n2132);
    or g560(n2427 ,n2271 ,n2131);
    or g561(n2426 ,n2270 ,n2130);
    or g562(n2425 ,n2269 ,n2129);
    or g563(n2424 ,n2268 ,n2128);
    or g564(n2423 ,n2267 ,n2172);
    or g565(n2422 ,n2266 ,n2127);
    or g566(n2421 ,n2265 ,n2126);
    or g567(n2420 ,n2264 ,n2125);
    or g568(n2419 ,n2263 ,n2124);
    or g569(n2418 ,n2262 ,n2123);
    or g570(n2417 ,n2261 ,n2122);
    or g571(n2416 ,n2260 ,n2121);
    or g572(n2415 ,n2259 ,n2171);
    or g573(n2414 ,n2257 ,n2119);
    or g574(n2413 ,n2258 ,n2120);
    or g575(n2412 ,n2256 ,n2118);
    or g576(n2411 ,n2255 ,n2117);
    or g577(n2410 ,n2254 ,n2116);
    or g578(n2409 ,n2253 ,n2115);
    or g579(n2408 ,n2252 ,n2114);
    or g580(n2407 ,n2251 ,n2332);
    or g581(n2406 ,n2250 ,n2062);
    or g582(n2405 ,n2280 ,n2061);
    or g583(n2404 ,n2249 ,n2060);
    or g584(n2403 ,n2248 ,n2059);
    or g585(n2402 ,n2335 ,n2058);
    or g586(n2401 ,n2246 ,n2057);
    or g587(n2400 ,n2245 ,n2056);
    or g588(n2399 ,n2244 ,n2170);
    or g589(n2398 ,n2242 ,n2112);
    or g590(n2397 ,n2243 ,n2113);
    or g591(n2396 ,n2241 ,n2111);
    or g592(n2395 ,n2240 ,n2110);
    or g593(n2394 ,n2239 ,n2109);
    or g594(n2393 ,n2238 ,n2108);
    or g595(n2392 ,n2237 ,n2107);
    or g596(n2391 ,n2236 ,n2169);
    or g597(n2390 ,n2235 ,n2106);
    or g598(n2389 ,n2234 ,n2105);
    or g599(n2388 ,n2233 ,n2104);
    or g600(n2387 ,n2232 ,n2103);
    or g601(n2386 ,n2231 ,n2102);
    or g602(n2385 ,n2229 ,n2100);
    or g603(n2384 ,n2230 ,n2101);
    or g604(n2383 ,n2228 ,n2168);
    or g605(n2382 ,n2227 ,n2099);
    or g606(n2381 ,n2226 ,n2098);
    or g607(n2380 ,n2225 ,n2097);
    or g608(n2379 ,n2224 ,n2096);
    or g609(n2378 ,n2223 ,n2095);
    or g610(n2377 ,n2222 ,n2094);
    or g611(n2376 ,n2221 ,n2093);
    or g612(n2375 ,n2220 ,n2167);
    or g613(n2374 ,n2219 ,n2092);
    or g614(n2373 ,n2218 ,n2091);
    or g615(n2372 ,n2217 ,n2090);
    or g616(n2371 ,n2216 ,n2089);
    or g617(n2370 ,n2215 ,n2088);
    or g618(n2369 ,n2214 ,n2087);
    or g619(n2368 ,n2213 ,n2086);
    or g620(n2367 ,n2212 ,n2247);
    or g621(n2366 ,n2211 ,n2085);
    or g622(n2365 ,n2210 ,n2084);
    or g623(n2364 ,n2209 ,n2083);
    or g624(n2363 ,n2207 ,n2082);
    or g625(n2362 ,n2208 ,n2081);
    or g626(n2361 ,n2206 ,n2080);
    or g627(n2360 ,n2205 ,n2079);
    or g628(n2359 ,n2204 ,n2329);
    or g629(n2358 ,n2203 ,n2078);
    or g630(n2357 ,n2202 ,n2077);
    or g631(n2356 ,n2201 ,n2076);
    or g632(n2355 ,n1478 ,n2316);
    or g633(n2354 ,n2200 ,n2075);
    or g634(n2353 ,n2199 ,n2074);
    or g635(n2352 ,n2198 ,n2073);
    or g636(n2351 ,n2197 ,n2072);
    or g637(n2350 ,n2196 ,n2330);
    or g638(n2349 ,n2195 ,n2071);
    or g639(n2348 ,n2194 ,n2070);
    or g640(n2347 ,n2193 ,n2069);
    or g641(n2346 ,n2192 ,n2068);
    or g642(n2345 ,n1485 ,n2315);
    or g643(n2344 ,n2191 ,n2067);
    or g644(n2343 ,n2190 ,n2066);
    or g645(n2342 ,n2189 ,n2065);
    or g646(n2341 ,n1482 ,n2048);
    or g647(n2340 ,n1481 ,n2314);
    or g648(n2339 ,n2188 ,n2331);
    or g649(n2338 ,n1479 ,n2317);
    or g650(n2337 ,n2187 ,n2064);
    or g651(n2336 ,n2186 ,n2063);
    nor g652(n2335 ,n434 ,n1879);
    nor g653(n2334 ,n290 ,n1908);
    nor g654(n2333 ,n289 ,n1908);
    nor g655(n2332 ,n497 ,n1878);
    nor g656(n2331 ,n497 ,n1908);
    nor g657(n2330 ,n497 ,n1906);
    nor g658(n2329 ,n497 ,n1902);
    nor g659(n2328 ,n444 ,n1911);
    nor g660(n2327 ,n455 ,n1911);
    nor g661(n2326 ,n470 ,n1911);
    nor g662(n2325 ,n451 ,n1910);
    nor g663(n2324 ,n484 ,n1910);
    nor g664(n2323 ,n493 ,n1910);
    nor g665(n2322 ,n456 ,n1910);
    nor g666(n2321 ,n458 ,n1910);
    nor g667(n2320 ,n467 ,n1910);
    nor g668(n2319 ,n462 ,n1910);
    nor g669(n2318 ,n473 ,n1910);
    nor g670(n2317 ,n471 ,n1910);
    nor g671(n2316 ,n466 ,n1910);
    nor g672(n2315 ,n454 ,n1910);
    nor g673(n2314 ,n460 ,n1910);
    nor g674(n2313 ,n671 ,n1909);
    nor g675(n2312 ,n393 ,n1909);
    nor g676(n2311 ,n408 ,n1909);
    nor g677(n2310 ,n536 ,n1909);
    nor g678(n2309 ,n630 ,n1909);
    nor g679(n2308 ,n697 ,n1881);
    nor g680(n2307 ,n635 ,n1881);
    nor g681(n2306 ,n332 ,n1881);
    nor g682(n2305 ,n689 ,n1881);
    nor g683(n2304 ,n640 ,n1881);
    nor g684(n2303 ,n608 ,n1881);
    nor g685(n2302 ,n568 ,n1881);
    nor g686(n2301 ,n593 ,n1881);
    nor g687(n2300 ,n331 ,n1883);
    nor g688(n2299 ,n538 ,n1883);
    nor g689(n2298 ,n428 ,n1883);
    nor g690(n2297 ,n380 ,n1883);
    nor g691(n2296 ,n352 ,n1883);
    nor g692(n2295 ,n655 ,n1883);
    nor g693(n2294 ,n441 ,n1883);
    nor g694(n2293 ,n574 ,n1883);
    nor g695(n2292 ,n628 ,n1885);
    nor g696(n2291 ,n383 ,n1885);
    nor g697(n2290 ,n578 ,n1885);
    nor g698(n2289 ,n690 ,n1885);
    nor g699(n2288 ,n615 ,n1885);
    nor g700(n2287 ,n351 ,n1885);
    nor g701(n2286 ,n558 ,n1885);
    nor g702(n2285 ,n580 ,n1885);
    nor g703(n2284 ,n329 ,n1887);
    nor g704(n2283 ,n410 ,n1887);
    nor g705(n2282 ,n319 ,n1887);
    nor g706(n2281 ,n415 ,n1887);
    nor g707(n2280 ,n379 ,n1879);
    nor g708(n2279 ,n409 ,n1887);
    nor g709(n2278 ,n346 ,n1887);
    nor g710(n2277 ,n321 ,n1887);
    nor g711(n2276 ,n318 ,n1887);
    nor g712(n2275 ,n406 ,n1889);
    nor g713(n2274 ,n663 ,n1889);
    nor g714(n2273 ,n657 ,n1889);
    nor g715(n2272 ,n335 ,n1889);
    nor g716(n2271 ,n605 ,n1889);
    nor g717(n2270 ,n670 ,n1889);
    nor g718(n2269 ,n327 ,n1889);
    nor g719(n2268 ,n362 ,n1889);
    nor g720(n2267 ,n582 ,n1895);
    nor g721(n2266 ,n439 ,n1895);
    nor g722(n2265 ,n560 ,n1895);
    nor g723(n2264 ,n609 ,n1895);
    nor g724(n2263 ,n339 ,n1895);
    nor g725(n2262 ,n579 ,n1895);
    nor g726(n2261 ,n585 ,n1895);
    nor g727(n2260 ,n653 ,n1895);
    nor g728(n2259 ,n624 ,n1891);
    nor g729(n2258 ,n665 ,n1891);
    nor g730(n2257 ,n540 ,n1891);
    nor g731(n2256 ,n396 ,n1891);
    nor g732(n2255 ,n324 ,n1891);
    nor g733(n2254 ,n334 ,n1891);
    nor g734(n2253 ,n427 ,n1891);
    nor g735(n2252 ,n694 ,n1891);
    nor g736(n2251 ,n562 ,n1879);
    nor g737(n2250 ,n357 ,n1879);
    nor g738(n2249 ,n433 ,n1879);
    nor g739(n2248 ,n375 ,n1879);
    nor g740(n2247 ,n497 ,n1900);
    nor g741(n2246 ,n399 ,n1879);
    nor g742(n2245 ,n641 ,n1879);
    nor g743(n2244 ,n599 ,n1893);
    nor g744(n2243 ,n696 ,n1893);
    nor g745(n2242 ,n418 ,n1893);
    nor g746(n2241 ,n389 ,n1893);
    nor g747(n2240 ,n422 ,n1893);
    nor g748(n2239 ,n348 ,n1893);
    nor g749(n2238 ,n432 ,n1893);
    nor g750(n2237 ,n692 ,n1893);
    nor g751(n2236 ,n645 ,n1905);
    nor g752(n2235 ,n386 ,n1905);
    nor g753(n2234 ,n364 ,n1905);
    nor g754(n2233 ,n576 ,n1905);
    nor g755(n2232 ,n438 ,n1905);
    nor g756(n2231 ,n551 ,n1905);
    nor g757(n2230 ,n367 ,n1905);
    nor g758(n2229 ,n384 ,n1905);
    nor g759(n2228 ,n682 ,n1897);
    nor g760(n2227 ,n344 ,n1897);
    nor g761(n2226 ,n548 ,n1897);
    nor g762(n2225 ,n440 ,n1897);
    nor g763(n2224 ,n606 ,n1897);
    nor g764(n2223 ,n337 ,n1897);
    nor g765(n2222 ,n636 ,n1897);
    nor g766(n2221 ,n350 ,n1897);
    nor g767(n2220 ,n584 ,n1899);
    nor g768(n2219 ,n354 ,n1899);
    nor g769(n2218 ,n398 ,n1899);
    nor g770(n2217 ,n591 ,n1899);
    nor g771(n2216 ,n349 ,n1899);
    nor g772(n2215 ,n442 ,n1899);
    nor g773(n2214 ,n649 ,n1899);
    nor g774(n2213 ,n661 ,n1899);
    nor g775(n2212 ,n559 ,n1901);
    nor g776(n2211 ,n650 ,n1901);
    nor g777(n2210 ,n631 ,n1901);
    nor g778(n2209 ,n426 ,n1901);
    nor g779(n2208 ,n589 ,n1901);
    nor g780(n2207 ,n382 ,n1901);
    nor g781(n2206 ,n674 ,n1901);
    nor g782(n2205 ,n683 ,n1901);
    nor g783(n2204 ,n413 ,n1903);
    nor g784(n2203 ,n372 ,n1903);
    nor g785(n2202 ,n412 ,n1903);
    nor g786(n2201 ,n361 ,n1903);
    nor g787(n2200 ,n684 ,n1903);
    nor g788(n2199 ,n676 ,n1903);
    nor g789(n2198 ,n668 ,n1903);
    nor g790(n2197 ,n403 ,n1903);
    nor g791(n2196 ,n400 ,n1907);
    nor g792(n2195 ,n627 ,n1907);
    nor g793(n2194 ,n687 ,n1907);
    nor g794(n2193 ,n660 ,n1907);
    nor g795(n2192 ,n378 ,n1907);
    nor g796(n2191 ,n537 ,n1907);
    nor g797(n2190 ,n647 ,n1907);
    nor g798(n2189 ,n654 ,n1907);
    nor g799(n2188 ,n385 ,n1909);
    nor g800(n2187 ,n358 ,n1909);
    nor g801(n2186 ,n643 ,n1909);
    or g802(n2185 ,n1203 ,n1808);
    or g803(n2184 ,n1183 ,n1807);
    or g804(n2183 ,n1179 ,n1810);
    or g805(n2182 ,n1173 ,n1805);
    or g806(n2181 ,n1163 ,n1809);
    or g807(n2180 ,n1161 ,n1804);
    or g808(n2179 ,n1141 ,n1811);
    or g809(n2178 ,n1184 ,n1812);
    nor g810(n2177 ,n497 ,n1880);
    nor g811(n2176 ,n497 ,n1882);
    nor g812(n2175 ,n497 ,n1884);
    nor g813(n2174 ,n497 ,n1886);
    nor g814(n2173 ,n497 ,n1888);
    nor g815(n2172 ,n497 ,n1894);
    nor g816(n2171 ,n497 ,n1890);
    nor g817(n2170 ,n497 ,n1892);
    nor g818(n2169 ,n497 ,n1904);
    nor g819(n2168 ,n497 ,n1896);
    nor g820(n2167 ,n497 ,n1898);
    or g821(n2165 ,n1837 ,n1923);
    nor g822(n2164 ,n288 ,n1908);
    nor g823(n2163 ,n495 ,n1908);
    nor g824(n2162 ,n287 ,n1880);
    nor g825(n2161 ,n496 ,n1880);
    nor g826(n2160 ,n289 ,n1880);
    nor g827(n2159 ,n290 ,n1880);
    nor g828(n2158 ,n494 ,n1880);
    nor g829(n2157 ,n288 ,n1880);
    nor g830(n2156 ,n495 ,n1880);
    nor g831(n2155 ,n287 ,n1882);
    nor g832(n2154 ,n496 ,n1882);
    nor g833(n2153 ,n289 ,n1882);
    nor g834(n2152 ,n290 ,n1882);
    nor g835(n2151 ,n494 ,n1882);
    nor g836(n2150 ,n288 ,n1882);
    nor g837(n2149 ,n495 ,n1882);
    nor g838(n2148 ,n287 ,n1884);
    nor g839(n2147 ,n496 ,n1884);
    nor g840(n2146 ,n289 ,n1884);
    nor g841(n2145 ,n290 ,n1884);
    nor g842(n2144 ,n494 ,n1884);
    nor g843(n2143 ,n288 ,n1884);
    nor g844(n2142 ,n495 ,n1884);
    nor g845(n2141 ,n287 ,n1886);
    nor g846(n2140 ,n496 ,n1886);
    nor g847(n2139 ,n289 ,n1886);
    nor g848(n2138 ,n290 ,n1886);
    nor g849(n2137 ,n494 ,n1886);
    nor g850(n2136 ,n288 ,n1886);
    nor g851(n2135 ,n495 ,n1886);
    nor g852(n2134 ,n287 ,n1888);
    nor g853(n2133 ,n496 ,n1888);
    nor g854(n2132 ,n289 ,n1888);
    nor g855(n2131 ,n290 ,n1888);
    nor g856(n2130 ,n494 ,n1888);
    nor g857(n2129 ,n288 ,n1888);
    nor g858(n2128 ,n495 ,n1888);
    nor g859(n2127 ,n287 ,n1894);
    nor g860(n2126 ,n496 ,n1894);
    nor g861(n2125 ,n289 ,n1894);
    nor g862(n2124 ,n290 ,n1894);
    nor g863(n2123 ,n494 ,n1894);
    nor g864(n2122 ,n288 ,n1894);
    nor g865(n2121 ,n495 ,n1894);
    nor g866(n2120 ,n287 ,n1890);
    nor g867(n2119 ,n496 ,n1890);
    nor g868(n2118 ,n289 ,n1890);
    nor g869(n2117 ,n290 ,n1890);
    nor g870(n2116 ,n494 ,n1890);
    nor g871(n2115 ,n288 ,n1890);
    nor g872(n2114 ,n495 ,n1890);
    nor g873(n2113 ,n287 ,n1892);
    nor g874(n2112 ,n496 ,n1892);
    nor g875(n2111 ,n289 ,n1892);
    nor g876(n2110 ,n290 ,n1892);
    nor g877(n2109 ,n494 ,n1892);
    nor g878(n2108 ,n288 ,n1892);
    nor g879(n2107 ,n495 ,n1892);
    nor g880(n2106 ,n287 ,n1904);
    nor g881(n2105 ,n496 ,n1904);
    nor g882(n2104 ,n289 ,n1904);
    nor g883(n2103 ,n290 ,n1904);
    nor g884(n2102 ,n494 ,n1904);
    nor g885(n2101 ,n288 ,n1904);
    nor g886(n2100 ,n495 ,n1904);
    nor g887(n2099 ,n287 ,n1896);
    nor g888(n2098 ,n496 ,n1896);
    nor g889(n2097 ,n289 ,n1896);
    nor g890(n2096 ,n290 ,n1896);
    nor g891(n2095 ,n494 ,n1896);
    nor g892(n2094 ,n288 ,n1896);
    nor g893(n2093 ,n495 ,n1896);
    nor g894(n2092 ,n287 ,n1898);
    nor g895(n2091 ,n496 ,n1898);
    nor g896(n2090 ,n289 ,n1898);
    nor g897(n2089 ,n290 ,n1898);
    nor g898(n2088 ,n494 ,n1898);
    nor g899(n2087 ,n288 ,n1898);
    nor g900(n2086 ,n495 ,n1898);
    nor g901(n2085 ,n287 ,n1900);
    nor g902(n2084 ,n496 ,n1900);
    nor g903(n2083 ,n289 ,n1900);
    nor g904(n2082 ,n290 ,n1900);
    nor g905(n2081 ,n494 ,n1900);
    nor g906(n2080 ,n288 ,n1900);
    nor g907(n2079 ,n495 ,n1900);
    nor g908(n2078 ,n287 ,n1902);
    nor g909(n2077 ,n496 ,n1902);
    nor g910(n2076 ,n289 ,n1902);
    nor g911(n2075 ,n290 ,n1902);
    nor g912(n2074 ,n494 ,n1902);
    nor g913(n2073 ,n288 ,n1902);
    nor g914(n2072 ,n495 ,n1902);
    nor g915(n2071 ,n287 ,n1906);
    nor g916(n2070 ,n496 ,n1906);
    nor g917(n2069 ,n289 ,n1906);
    nor g918(n2068 ,n290 ,n1906);
    nor g919(n2067 ,n494 ,n1906);
    nor g920(n2066 ,n288 ,n1906);
    nor g921(n2065 ,n495 ,n1906);
    nor g922(n2064 ,n287 ,n1908);
    nor g923(n2063 ,n496 ,n1908);
    nor g924(n2062 ,n287 ,n1878);
    nor g925(n2061 ,n496 ,n1878);
    nor g926(n2060 ,n289 ,n1878);
    nor g927(n2059 ,n290 ,n1878);
    nor g928(n2058 ,n494 ,n1878);
    nor g929(n2057 ,n288 ,n1878);
    nor g930(n2056 ,n495 ,n1878);
    nor g931(n2055 ,n494 ,n1908);
    nor g932(n2054 ,n281 ,n1820);
    nor g933(n2053 ,n286 ,n1821);
    nor g934(n2052 ,n286 ,n1822);
    nor g935(n2051 ,n284 ,n1823);
    nor g936(n2050 ,n286 ,n1824);
    nor g937(n2049 ,n285 ,n1825);
    nor g938(n2048 ,n20[0] ,n1910);
    or g939(n2047 ,n1871 ,n1855);
    or g940(n2046 ,n1965 ,n1987);
    or g941(n2045 ,n1986 ,n1960);
    or g942(n2044 ,n1984 ,n1962);
    or g943(n2043 ,n1955 ,n1954);
    or g944(n2042 ,n1952 ,n1716);
    or g945(n2041 ,n1951 ,n1950);
    or g946(n2040 ,n1864 ,n1918);
    or g947(n2039 ,n1964 ,n1947);
    or g948(n2038 ,n1967 ,n1946);
    or g949(n2037 ,n1969 ,n1944);
    or g950(n2036 ,n1989 ,n1942);
    or g951(n2035 ,n1940 ,n1939);
    or g952(n2034 ,n1938 ,n1714);
    or g953(n2033 ,n1937 ,n1912);
    or g954(n2032 ,n1934 ,n1936);
    or g955(n2031 ,n1933 ,n1953);
    or g956(n2030 ,n1856 ,n1931);
    or g957(n2029 ,n1935 ,n1948);
    or g958(n2028 ,n1741 ,n1806);
    or g959(n2027 ,n1858 ,n1715);
    or g960(n2026 ,n1861 ,n1927);
    or g961(n2025 ,n1845 ,n1836);
    or g962(n2024 ,n1925 ,n1924);
    or g963(n2023 ,n1834 ,n1835);
    or g964(n2022 ,n1840 ,n1838);
    or g965(n2021 ,n1739 ,n1975);
    or g966(n2020 ,n1919 ,n1844);
    or g967(n2019 ,n1846 ,n1847);
    or g968(n2018 ,n1917 ,n1848);
    or g969(n2017 ,n1915 ,n1849);
    or g970(n2016 ,n1850 ,n1851);
    or g971(n2015 ,n1958 ,n1922);
    or g972(n2014 ,n1913 ,n1945);
    or g973(n2013 ,n1875 ,n1711);
    or g974(n2012 ,n1862 ,n1865);
    or g975(n2011 ,n1976 ,n1985);
    or g976(n2010 ,n1740 ,n1974);
    or g977(n2009 ,n1831 ,n1977);
    or g978(n2008 ,n1979 ,n1916);
    or g979(n2007 ,n1981 ,n1978);
    or g980(n2006 ,n1982 ,n1712);
    or g981(n2005 ,n1961 ,n1966);
    or g982(n2004 ,n1957 ,n1959);
    or g983(n2003 ,n1841 ,n1863);
    or g984(n2002 ,n1876 ,n1968);
    or g985(n2001 ,n1970 ,n1713);
    or g986(n2000 ,n1972 ,n1873);
    or g987(n1999 ,n1857 ,n1973);
    or g988(n1998 ,n1870 ,n1949);
    or g989(n1997 ,n1869 ,n1929);
    or g990(n1996 ,n1867 ,n1709);
    or g991(n1995 ,n1854 ,n1866);
    or g992(n1994 ,n1842 ,n1980);
    or g993(n1993 ,n1988 ,n1843);
    or g994(n1992 ,n1932 ,n1860);
    or g995(n1991 ,n1920 ,n1710);
    or g996(n1990 ,n1928 ,n1859);
    nor g997(n1989 ,n644 ,n1784);
    nor g998(n1988 ,n695 ,n1784);
    nor g999(n1987 ,n360 ,n1789);
    nor g1000(n1986 ,n336 ,n1797);
    nor g1001(n1985 ,n419 ,n1785);
    nor g1002(n1984 ,n430 ,n1787);
    nor g1003(n1983 ,n387 ,n1788);
    nor g1004(n1982 ,n622 ,n1791);
    nor g1005(n1981 ,n326 ,n1797);
    nor g1006(n1980 ,n667 ,n1798);
    nor g1007(n1979 ,n681 ,n1784);
    nor g1008(n1978 ,n392 ,n1798);
    nor g1009(n1977 ,n617 ,n1786);
    nor g1010(n1976 ,n363 ,n1795);
    nor g1011(n1975 ,n463 ,n1803);
    nor g1012(n1974 ,n490 ,n1803);
    nor g1013(n1973 ,n417 ,n1786);
    nor g1014(n1972 ,n435 ,n1790);
    nor g1015(n1971 ,n625 ,n1792);
    nor g1016(n1970 ,n394 ,n1791);
    nor g1017(n1969 ,n338 ,n1797);
    nor g1018(n1968 ,n563 ,n1796);
    nor g1019(n1967 ,n620 ,n1787);
    nor g1020(n1966 ,n595 ,n1794);
    nor g1021(n1965 ,n586 ,n1784);
    nor g1022(n1964 ,n570 ,n1795);
    nor g1023(n1963 ,n353 ,n1788);
    nor g1024(n1962 ,n322 ,n1786);
    nor g1025(n1961 ,n588 ,n1790);
    nor g1026(n1960 ,n677 ,n1798);
    nor g1027(n1959 ,n342 ,n1785);
    nor g1028(n1958 ,n679 ,n1793);
    nor g1029(n1957 ,n391 ,n1795);
    nor g1030(n1956 ,n600 ,n1792);
    nor g1031(n1955 ,n632 ,n1793);
    nor g1032(n1954 ,n601 ,n1796);
    nor g1033(n1953 ,n368 ,n1786);
    nor g1034(n1952 ,n592 ,n1791);
    nor g1035(n1951 ,n637 ,n1790);
    nor g1036(n1950 ,n646 ,n1794);
    nor g1037(n1949 ,n374 ,n1798);
    nor g1038(n1948 ,n341 ,n1796);
    nor g1039(n1947 ,n597 ,n1785);
    nor g1040(n1946 ,n583 ,n1786);
    nor g1041(n1945 ,n425 ,n1796);
    nor g1042(n1944 ,n633 ,n1798);
    nor g1043(n1943 ,n602 ,n1788);
    nor g1044(n1942 ,n369 ,n1789);
    nor g1045(n1941 ,n691 ,n1792);
    nor g1046(n1940 ,n648 ,n1793);
    nor g1047(n1939 ,n539 ,n1796);
    nor g1048(n1938 ,n544 ,n1791);
    nor g1049(n1937 ,n365 ,n1790);
    nor g1050(n1936 ,n552 ,n1785);
    nor g1051(n1935 ,n557 ,n1793);
    nor g1052(n1934 ,n565 ,n1795);
    nor g1053(n1933 ,n554 ,n1787);
    nor g1054(n1932 ,n404 ,n1797);
    nor g1055(n1931 ,n581 ,n1789);
    nor g1056(n1930 ,n373 ,n1792);
    nor g1057(n1929 ,n561 ,n1789);
    nor g1058(n1928 ,n405 ,n1793);
    nor g1059(n1927 ,n693 ,n1794);
    nor g1060(n1926 ,n366 ,n1788);
    nor g1061(n1925 ,n541 ,n1787);
    nor g1062(n1924 ,n673 ,n1786);
    nor g1063(n1923 ,n611 ,n1789);
    nor g1064(n1922 ,n685 ,n1796);
    nor g1065(n1921 ,n395 ,n1788);
    nor g1066(n1920 ,n345 ,n1791);
    nor g1067(n1919 ,n370 ,n1790);
    nor g1068(n1918 ,n443 ,n1785);
    nor g1069(n1917 ,n555 ,n1787);
    nor g1070(n1916 ,n377 ,n1789);
    nor g1071(n1915 ,n623 ,n1797);
    nor g1072(n1914 ,n414 ,n1792);
    nor g1073(n1913 ,n381 ,n1793);
    nor g1074(n1912 ,n437 ,n1794);
    not g1075(n1908 ,n1909);
    not g1076(n1906 ,n1907);
    not g1077(n1904 ,n1905);
    not g1078(n1902 ,n1903);
    not g1079(n1900 ,n1901);
    not g1080(n1898 ,n1899);
    not g1081(n1896 ,n1897);
    not g1082(n1894 ,n1895);
    not g1083(n1892 ,n1893);
    not g1084(n1890 ,n1891);
    not g1085(n1888 ,n1889);
    not g1086(n1886 ,n1887);
    not g1087(n1884 ,n1885);
    not g1088(n1882 ,n1883);
    not g1089(n1880 ,n1881);
    not g1090(n1878 ,n1879);
    nor g1091(n1877 ,n416 ,n1783);
    nor g1092(n1876 ,n546 ,n1793);
    nor g1093(n1875 ,n634 ,n1791);
    nor g1094(n1874 ,n355 ,n1788);
    nor g1095(n1873 ,n598 ,n1794);
    nor g1096(n1872 ,n553 ,n1788);
    nor g1097(n1871 ,n388 ,n1795);
    nor g1098(n1870 ,n669 ,n1797);
    nor g1099(n1869 ,n662 ,n1784);
    nor g1100(n1868 ,n658 ,n1792);
    nor g1101(n1867 ,n619 ,n1791);
    nor g1102(n1866 ,n621 ,n1794);
    nor g1103(n1865 ,n666 ,n1794);
    nor g1104(n1864 ,n397 ,n1795);
    nor g1105(n1863 ,n614 ,n1786);
    nor g1106(n1862 ,n664 ,n1790);
    nor g1107(n1861 ,n347 ,n1790);
    nor g1108(n1860 ,n569 ,n1798);
    nor g1109(n1859 ,n429 ,n1796);
    nor g1110(n1858 ,n612 ,n1791);
    nor g1111(n1857 ,n577 ,n1787);
    nor g1112(n1856 ,n402 ,n1784);
    nor g1113(n1855 ,n340 ,n1785);
    nor g1114(n1854 ,n356 ,n1790);
    nor g1115(n1853 ,n564 ,n1792);
    nor g1116(n1852 ,n680 ,n1788);
    nor g1117(n1851 ,n596 ,n1789);
    nor g1118(n1850 ,n567 ,n1784);
    nor g1119(n1849 ,n371 ,n1798);
    nor g1120(n1848 ,n688 ,n1786);
    nor g1121(n1847 ,n571 ,n1785);
    nor g1122(n1846 ,n436 ,n1795);
    nor g1123(n1845 ,n343 ,n1795);
    nor g1124(n1844 ,n610 ,n1794);
    nor g1125(n1843 ,n607 ,n1789);
    nor g1126(n1842 ,n411 ,n1797);
    nor g1127(n1841 ,n652 ,n1787);
    nor g1128(n1840 ,n659 ,n1793);
    nor g1129(n1839 ,n547 ,n1792);
    nor g1130(n1838 ,n587 ,n1796);
    nor g1131(n1837 ,n616 ,n1784);
    nor g1132(n1836 ,n572 ,n1785);
    nor g1133(n1835 ,n613 ,n1798);
    nor g1134(n1834 ,n333 ,n1797);
    nor g1135(n1833 ,n401 ,n1783);
    nor g1136(n1832 ,n421 ,n1783);
    nor g1137(n1831 ,n651 ,n1787);
    nor g1138(n1830 ,n594 ,n1783);
    nor g1139(n1829 ,n325 ,n1783);
    nor g1140(n1828 ,n323 ,n1783);
    nor g1141(n1827 ,n556 ,n1783);
    nor g1142(n1826 ,n407 ,n1783);
    nor g1143(n1825 ,n1754 ,n1762);
    nor g1144(n1824 ,n892 ,n1753);
    nor g1145(n1823 ,n1743 ,n1761);
    nor g1146(n1822 ,n1752 ,n1760);
    nor g1147(n1821 ,n1742 ,n1759);
    nor g1148(n1820 ,n1738 ,n1758);
    nor g1149(n1819 ,n282 ,n1777);
    nor g1150(n1818 ,n282 ,n1773);
    nor g1151(n1817 ,n281 ,n1772);
    nor g1152(n1816 ,n282 ,n1771);
    nor g1153(n1815 ,n280 ,n1775);
    nor g1154(n1814 ,n284 ,n1767);
    nor g1155(n1813 ,n282 ,n1781);
    or g1156(n1812 ,n801 ,n1751);
    or g1157(n1811 ,n803 ,n1750);
    or g1158(n1810 ,n800 ,n1745);
    or g1159(n1809 ,n802 ,n1749);
    or g1160(n1808 ,n806 ,n1744);
    or g1161(n1807 ,n765 ,n1746);
    nor g1162(n1806 ,n18[0] ,n1803);
    or g1163(n1805 ,n805 ,n1747);
    or g1164(n1804 ,n798 ,n1748);
    or g1165(n1911 ,n1036 ,n1782);
    or g1166(n1910 ,n286 ,n1763);
    nor g1167(n1909 ,n748 ,n1800);
    nor g1168(n1907 ,n748 ,n1801);
    nor g1169(n1905 ,n717 ,n1800);
    nor g1170(n1903 ,n715 ,n1800);
    nor g1171(n1901 ,n715 ,n1801);
    nor g1172(n1899 ,n713 ,n1800);
    nor g1173(n1897 ,n713 ,n1801);
    nor g1174(n1895 ,n715 ,n1799);
    nor g1175(n1893 ,n717 ,n1801);
    nor g1176(n1891 ,n748 ,n1802);
    nor g1177(n1889 ,n715 ,n1802);
    nor g1178(n1887 ,n713 ,n1799);
    nor g1179(n1885 ,n713 ,n1802);
    nor g1180(n1883 ,n717 ,n1799);
    nor g1181(n1881 ,n717 ,n1802);
    nor g1182(n1879 ,n748 ,n1799);
    not g1183(n1783 ,n1782);
    xnor g1184(n1781 ,n1322 ,n19[0]);
    or g1185(n1780 ,n759 ,n1670);
    or g1186(n1779 ,n1720 ,n1719);
    or g1187(n1778 ,n1722 ,n1721);
    nor g1188(n1777 ,n1669 ,n1723);
    or g1189(n1776 ,n1701 ,n1663);
    nor g1190(n1775 ,n1705 ,n1708);
    or g1191(n1774 ,n1717 ,n1735);
    nor g1192(n1773 ,n1702 ,n1698);
    nor g1193(n1772 ,n1703 ,n1706);
    nor g1194(n1771 ,n1704 ,n1707);
    or g1195(n1770 ,n845 ,n1725);
    or g1196(n1769 ,n848 ,n1724);
    or g1197(n1768 ,n857 ,n1726);
    nor g1198(n1767 ,n1506 ,n1666);
    nor g1199(n1766 ,n283 ,n1612);
    nor g1200(n1765 ,n280 ,n1613);
    or g1201(n1764 ,n1495 ,n1530);
    or g1202(n1763 ,n894 ,n1557);
    nor g1203(n1762 ,n729 ,n1626);
    nor g1204(n1761 ,n794 ,n1626);
    nor g1205(n1760 ,n707 ,n1729);
    nor g1206(n1759 ,n762 ,n1729);
    nor g1207(n1758 ,n785 ,n1729);
    or g1208(n1757 ,n1492 ,n1624);
    or g1209(n1756 ,n1494 ,n1570);
    or g1210(n1755 ,n1491 ,n1718);
    nor g1211(n1754 ,n498 ,n1627);
    nor g1212(n1753 ,n499 ,n1627);
    nor g1213(n1752 ,n299 ,n1728);
    or g1214(n1751 ,n1672 ,n1671);
    or g1215(n1750 ,n1676 ,n1675);
    or g1216(n1749 ,n1682 ,n1680);
    or g1217(n1748 ,n1684 ,n1683);
    or g1218(n1747 ,n1687 ,n1686);
    or g1219(n1746 ,n1677 ,n1690);
    or g1220(n1745 ,n1691 ,n1681);
    or g1221(n1744 ,n1693 ,n1692);
    nor g1222(n1743 ,n500 ,n1627);
    nor g1223(n1742 ,n307 ,n1728);
    nor g1224(n1741 ,n512 ,n1734);
    nor g1225(n1740 ,n317 ,n1734);
    nor g1226(n1739 ,n523 ,n1734);
    nor g1227(n1738 ,n308 ,n1728);
    or g1228(n1803 ,n881 ,n1665);
    or g1229(n1802 ,n505 ,n1736);
    or g1230(n1801 ,n38[3] ,n1736);
    or g1231(n1800 ,n38[3] ,n1737);
    or g1232(n1799 ,n505 ,n1737);
    or g1233(n1798 ,n721 ,n1730);
    or g1234(n1797 ,n721 ,n1732);
    or g1235(n1796 ,n721 ,n1733);
    or g1236(n1795 ,n749 ,n1730);
    or g1237(n1794 ,n716 ,n1733);
    or g1238(n1793 ,n721 ,n1731);
    or g1239(n1792 ,n719 ,n1731);
    or g1240(n1791 ,n749 ,n1732);
    or g1241(n1790 ,n716 ,n1731);
    or g1242(n1789 ,n719 ,n1730);
    or g1243(n1788 ,n749 ,n1733);
    or g1244(n1787 ,n716 ,n1732);
    or g1245(n1786 ,n716 ,n1730);
    or g1246(n1785 ,n719 ,n1733);
    or g1247(n1784 ,n719 ,n1732);
    nor g1248(n1782 ,n749 ,n1731);
    not g1249(n1736 ,n1735);
    not g1250(n1728 ,n1729);
    or g1251(n1727 ,n1207 ,n1205);
    nor g1252(n1726 ,n477 ,n1326);
    nor g1253(n1725 ,n450 ,n1326);
    nor g1254(n1724 ,n472 ,n1326);
    nor g1255(n1723 ,n524 ,n1331);
    nor g1256(n1722 ,n514 ,n1327);
    nor g1257(n1721 ,n475 ,n1515);
    nor g1258(n1720 ,n310 ,n1327);
    nor g1259(n1719 ,n481 ,n1515);
    or g1260(n1718 ,n854 ,n1498);
    nor g1261(n1717 ,n513 ,n1325);
    nor g1262(n1716 ,n543 ,n1324);
    nor g1263(n1715 ,n573 ,n1324);
    nor g1264(n1714 ,n545 ,n1324);
    nor g1265(n1713 ,n590 ,n1324);
    nor g1266(n1712 ,n424 ,n1324);
    nor g1267(n1711 ,n549 ,n1324);
    nor g1268(n1710 ,n604 ,n1324);
    nor g1269(n1709 ,n603 ,n1324);
    nor g1270(n1708 ,n529 ,n1322);
    nor g1271(n1707 ,n532 ,n1322);
    nor g1272(n1706 ,n525 ,n1322);
    nor g1273(n1705 ,n447 ,n1323);
    nor g1274(n1704 ,n485 ,n1323);
    nor g1275(n1703 ,n483 ,n1323);
    nor g1276(n1702 ,n474 ,n1323);
    nor g1277(n1701 ,n510 ,n1327);
    or g1278(n1700 ,n1452 ,n1215);
    or g1279(n1699 ,n1450 ,n1216);
    nor g1280(n1698 ,n511 ,n1322);
    nor g1281(n1697 ,n504 ,n1325);
    nor g1282(n1696 ,n506 ,n1325);
    nor g1283(n1695 ,n505 ,n1325);
    or g1284(n1694 ,n1197 ,n1204);
    or g1285(n1693 ,n1181 ,n1190);
    or g1286(n1692 ,n1200 ,n1189);
    or g1287(n1691 ,n1196 ,n1199);
    or g1288(n1690 ,n1191 ,n1188);
    or g1289(n1689 ,n1175 ,n1174);
    or g1290(n1688 ,n1170 ,n1166);
    or g1291(n1687 ,n1171 ,n1169);
    or g1292(n1686 ,n1168 ,n1167);
    or g1293(n1685 ,n1165 ,n1164);
    or g1294(n1684 ,n1157 ,n1155);
    or g1295(n1683 ,n1151 ,n1147);
    or g1296(n1682 ,n1149 ,n1145);
    or g1297(n1681 ,n1192 ,n1182);
    or g1298(n1680 ,n1143 ,n1198);
    or g1299(n1679 ,n1202 ,n1187);
    or g1300(n1678 ,n1140 ,n1195);
    or g1301(n1677 ,n1193 ,n1177);
    or g1302(n1676 ,n1172 ,n1201);
    or g1303(n1675 ,n1144 ,n1180);
    or g1304(n1674 ,n1178 ,n1176);
    or g1305(n1673 ,n1455 ,n1220);
    or g1306(n1672 ,n1210 ,n1206);
    or g1307(n1671 ,n1208 ,n1185);
    nor g1308(n1670 ,n931 ,n1325);
    nor g1309(n1669 ,n498 ,n1330);
    or g1310(n1668 ,n1445 ,n1217);
    or g1311(n1667 ,n1456 ,n1214);
    nor g1312(n1666 ,n17[2] ,n1186);
    or g1313(n1665 ,n892 ,n1333);
    or g1314(n1664 ,n1441 ,n1218);
    nor g1315(n1663 ,n41[0] ,n1515);
    or g1316(n1662 ,n1457 ,n1219);
    or g1317(n1661 ,n1459 ,n1513);
    nor g1318(n1660 ,n285 ,n1321);
    nor g1319(n1659 ,n284 ,n1162);
    nor g1320(n1658 ,n283 ,n1160);
    nor g1321(n1657 ,n280 ,n1159);
    nor g1322(n1656 ,n283 ,n1158);
    nor g1323(n1655 ,n281 ,n1156);
    nor g1324(n1654 ,n281 ,n1154);
    nor g1325(n1653 ,n280 ,n1153);
    nor g1326(n1652 ,n285 ,n1152);
    nor g1327(n1651 ,n284 ,n1150);
    nor g1328(n1650 ,n285 ,n1148);
    nor g1329(n1649 ,n280 ,n1146);
    or g1330(n1648 ,n1476 ,n1342);
    or g1331(n1647 ,n1475 ,n1341);
    or g1332(n1646 ,n1474 ,n1514);
    or g1333(n1645 ,n1472 ,n1340);
    or g1334(n1644 ,n1471 ,n1339);
    or g1335(n1643 ,n1435 ,n1338);
    or g1336(n1642 ,n1470 ,n1252);
    or g1337(n1641 ,n1469 ,n1337);
    or g1338(n1640 ,n1468 ,n1336);
    or g1339(n1639 ,n1467 ,n1284);
    or g1340(n1638 ,n1466 ,n1306);
    or g1341(n1637 ,n1414 ,n1334);
    or g1342(n1636 ,n1465 ,n1318);
    or g1343(n1635 ,n1464 ,n1346);
    or g1344(n1634 ,n1439 ,n1493);
    or g1345(n1633 ,n1463 ,n1507);
    or g1346(n1632 ,n1462 ,n1508);
    or g1347(n1631 ,n1442 ,n1509);
    or g1348(n1630 ,n1461 ,n1213);
    or g1349(n1629 ,n1446 ,n1510);
    or g1350(n1628 ,n1448 ,n1512);
    or g1351(n1737 ,n513 ,n1328);
    nor g1352(n1735 ,n38[0] ,n1328);
    or g1353(n1734 ,n278 ,n1332);
    or g1354(n1733 ,n59[0] ,n1516);
    or g1355(n1732 ,n501 ,n1329);
    or g1356(n1731 ,n501 ,n1516);
    or g1357(n1730 ,n59[0] ,n1329);
    nor g1358(n1729 ,n1194 ,n1044);
    not g1359(n1627 ,n1626);
    or g1360(n1625 ,n1390 ,n1335);
    or g1361(n1624 ,n853 ,n1347);
    or g1362(n1623 ,n1460 ,n1511);
    or g1363(n1622 ,n1447 ,n1262);
    or g1364(n1621 ,n1402 ,n1286);
    or g1365(n1620 ,n1356 ,n1232);
    or g1366(n1619 ,n1458 ,n1320);
    or g1367(n1618 ,n776 ,n1505);
    or g1368(n1617 ,n777 ,n1504);
    or g1369(n1616 ,n799 ,n1503);
    or g1370(n1615 ,n1454 ,n1221);
    or g1371(n1614 ,n1477 ,n1343);
    nor g1372(n1613 ,n1142 ,n1502);
    nor g1373(n1612 ,n1344 ,n1501);
    or g1374(n1611 ,n1431 ,n1317);
    or g1375(n1610 ,n1430 ,n1316);
    or g1376(n1609 ,n1429 ,n1315);
    or g1377(n1608 ,n1428 ,n1314);
    or g1378(n1607 ,n1427 ,n1312);
    or g1379(n1606 ,n1426 ,n1311);
    or g1380(n1605 ,n1425 ,n1310);
    or g1381(n1604 ,n1424 ,n1309);
    or g1382(n1603 ,n1423 ,n1308);
    or g1383(n1602 ,n1422 ,n1307);
    or g1384(n1601 ,n1421 ,n1304);
    or g1385(n1600 ,n1420 ,n1303);
    or g1386(n1599 ,n1419 ,n1302);
    or g1387(n1598 ,n1418 ,n1301);
    or g1388(n1597 ,n1417 ,n1300);
    or g1389(n1596 ,n1416 ,n1299);
    or g1390(n1595 ,n1415 ,n1298);
    or g1391(n1594 ,n1453 ,n1297);
    or g1392(n1593 ,n1413 ,n1296);
    or g1393(n1592 ,n1412 ,n1295);
    or g1394(n1591 ,n1410 ,n1294);
    or g1395(n1590 ,n1409 ,n1293);
    or g1396(n1589 ,n1408 ,n1292);
    or g1397(n1588 ,n1432 ,n1291);
    or g1398(n1587 ,n1406 ,n1290);
    or g1399(n1586 ,n1405 ,n1313);
    or g1400(n1585 ,n1433 ,n1289);
    or g1401(n1584 ,n1404 ,n1288);
    or g1402(n1583 ,n1403 ,n1287);
    or g1403(n1582 ,n1411 ,n1235);
    or g1404(n1581 ,n1401 ,n1285);
    or g1405(n1580 ,n1400 ,n1283);
    or g1406(n1579 ,n1399 ,n1282);
    or g1407(n1578 ,n1398 ,n1281);
    or g1408(n1577 ,n1397 ,n1280);
    or g1409(n1576 ,n1396 ,n1279);
    or g1410(n1575 ,n1395 ,n1278);
    or g1411(n1574 ,n1394 ,n1277);
    or g1412(n1573 ,n1393 ,n1276);
    or g1413(n1572 ,n1392 ,n1275);
    or g1414(n1571 ,n1437 ,n1274);
    or g1415(n1570 ,n852 ,n1496);
    or g1416(n1569 ,n1438 ,n1273);
    or g1417(n1568 ,n1391 ,n1319);
    or g1418(n1567 ,n1440 ,n1272);
    or g1419(n1566 ,n1389 ,n1271);
    or g1420(n1565 ,n1388 ,n1270);
    or g1421(n1564 ,n1387 ,n1269);
    or g1422(n1563 ,n1386 ,n1268);
    or g1423(n1562 ,n1385 ,n1267);
    or g1424(n1561 ,n1444 ,n1266);
    or g1425(n1560 ,n1384 ,n1265);
    or g1426(n1559 ,n1383 ,n1264);
    or g1427(n1558 ,n1382 ,n1263);
    nor g1428(n1557 ,n767 ,n1209);
    or g1429(n1556 ,n1381 ,n1261);
    or g1430(n1555 ,n1380 ,n1305);
    or g1431(n1554 ,n1379 ,n1260);
    or g1432(n1553 ,n1378 ,n1259);
    or g1433(n1552 ,n1377 ,n1258);
    or g1434(n1551 ,n1375 ,n1257);
    or g1435(n1550 ,n1436 ,n1256);
    or g1436(n1549 ,n1374 ,n1255);
    or g1437(n1548 ,n1373 ,n1254);
    or g1438(n1547 ,n1372 ,n1253);
    or g1439(n1546 ,n1371 ,n1251);
    or g1440(n1545 ,n1370 ,n1250);
    or g1441(n1544 ,n1369 ,n1249);
    or g1442(n1543 ,n1368 ,n1248);
    or g1443(n1542 ,n1367 ,n1247);
    or g1444(n1541 ,n1451 ,n1246);
    or g1445(n1540 ,n1366 ,n1245);
    or g1446(n1539 ,n1434 ,n1244);
    or g1447(n1538 ,n1365 ,n1243);
    or g1448(n1537 ,n1364 ,n1242);
    or g1449(n1536 ,n1363 ,n1241);
    or g1450(n1535 ,n1376 ,n1240);
    or g1451(n1534 ,n1362 ,n1239);
    or g1452(n1533 ,n1361 ,n1238);
    or g1453(n1532 ,n1360 ,n1237);
    or g1454(n1531 ,n1407 ,n1236);
    or g1455(n1530 ,n855 ,n1497);
    or g1456(n1529 ,n1358 ,n1234);
    or g1457(n1528 ,n1357 ,n1233);
    or g1458(n1527 ,n1355 ,n1231);
    or g1459(n1526 ,n1354 ,n1230);
    or g1460(n1525 ,n1443 ,n1229);
    or g1461(n1524 ,n1353 ,n1228);
    or g1462(n1523 ,n1499 ,n1211);
    or g1463(n1522 ,n1449 ,n1227);
    or g1464(n1521 ,n1352 ,n1226);
    or g1465(n1520 ,n1351 ,n1225);
    or g1466(n1519 ,n1350 ,n1224);
    or g1467(n1518 ,n1473 ,n1223);
    or g1468(n1517 ,n1359 ,n1222);
    nor g1469(n1626 ,n1212 ,n933);
    nor g1470(n1514 ,n291 ,n1019);
    nor g1471(n1513 ,n298 ,n1009);
    nor g1472(n1512 ,n296 ,n1009);
    nor g1473(n1511 ,n292 ,n1009);
    nor g1474(n1510 ,n294 ,n1009);
    nor g1475(n1509 ,n297 ,n1009);
    nor g1476(n1508 ,n291 ,n1009);
    nor g1477(n1507 ,n295 ,n1009);
    nor g1478(n1506 ,n517 ,n1046);
    nor g1479(n1505 ,n487 ,n1042);
    nor g1480(n1504 ,n453 ,n1042);
    nor g1481(n1503 ,n448 ,n1042);
    nor g1482(n1502 ,n530 ,n1044);
    nor g1483(n1501 ,n533 ,n1048);
    nor g1484(n1500 ,n515 ,n1039);
    nor g1485(n1499 ,n534 ,n1038);
    nor g1486(n1498 ,n528 ,n1038);
    nor g1487(n1497 ,n519 ,n1038);
    nor g1488(n1496 ,n527 ,n1038);
    nor g1489(n1495 ,n486 ,n1036);
    nor g1490(n1494 ,n445 ,n1036);
    nor g1491(n1493 ,n298 ,n1011);
    nor g1492(n1492 ,n469 ,n1036);
    nor g1493(n1491 ,n492 ,n1036);
    nor g1494(n1490 ,n686 ,n1035);
    nor g1495(n1489 ,n629 ,n1035);
    nor g1496(n1488 ,n656 ,n1035);
    nor g1497(n1487 ,n638 ,n1035);
    nor g1498(n1486 ,n642 ,n1035);
    nor g1499(n1485 ,n566 ,n1035);
    nor g1500(n1484 ,n423 ,n1035);
    nor g1501(n1483 ,n542 ,n1035);
    nor g1502(n1482 ,n522 ,n1035);
    nor g1503(n1481 ,n359 ,n1035);
    nor g1504(n1480 ,n431 ,n1035);
    nor g1505(n1479 ,n550 ,n1035);
    nor g1506(n1478 ,n618 ,n1035);
    nor g1507(n1477 ,n546 ,n1014);
    nor g1508(n1476 ,n679 ,n1014);
    nor g1509(n1475 ,n646 ,n1020);
    nor g1510(n1474 ,n437 ,n1020);
    nor g1511(n1473 ,n381 ,n1014);
    nor g1512(n1472 ,n693 ,n1020);
    nor g1513(n1471 ,n610 ,n1020);
    nor g1514(n1470 ,n595 ,n1020);
    nor g1515(n1469 ,n598 ,n1020);
    nor g1516(n1468 ,n621 ,n1020);
    nor g1517(n1467 ,n365 ,n1012);
    nor g1518(n1466 ,n347 ,n1012);
    nor g1519(n1465 ,n664 ,n1012);
    nor g1520(n1464 ,n588 ,n1012);
    nor g1521(n1463 ,n353 ,n1010);
    nor g1522(n1462 ,n395 ,n1010);
    nor g1523(n1461 ,n680 ,n1010);
    nor g1524(n1460 ,n387 ,n1010);
    nor g1525(n1459 ,n355 ,n1010);
    nor g1526(n1458 ,n435 ,n1012);
    nor g1527(n1457 ,n416 ,n1004);
    nor g1528(n1456 ,n323 ,n1004);
    nor g1529(n1455 ,n407 ,n1004);
    nor g1530(n1454 ,n401 ,n1004);
    nor g1531(n1453 ,n569 ,n1030);
    nor g1532(n1452 ,n556 ,n1004);
    nor g1533(n1451 ,n342 ,n1008);
    nor g1534(n1450 ,n421 ,n1004);
    nor g1535(n1449 ,n632 ,n1014);
    nor g1536(n1448 ,n553 ,n1010);
    nor g1537(n1447 ,n391 ,n1006);
    nor g1538(n1446 ,n602 ,n1010);
    nor g1539(n1445 ,n325 ,n1004);
    nor g1540(n1444 ,n565 ,n1006);
    nor g1541(n1443 ,n563 ,n1028);
    nor g1542(n1442 ,n366 ,n1010);
    nor g1543(n1441 ,n594 ,n1004);
    nor g1544(n1440 ,n555 ,n1034);
    nor g1545(n1439 ,n356 ,n1012);
    nor g1546(n1438 ,n554 ,n1034);
    nor g1547(n1437 ,n620 ,n1034);
    nor g1548(n1436 ,n634 ,n1018);
    nor g1549(n1435 ,n666 ,n1020);
    nor g1550(n1434 ,n443 ,n1008);
    nor g1551(n1433 ,n333 ,n1016);
    nor g1552(n1432 ,n667 ,n1030);
    nor g1553(n1431 ,n369 ,n1022);
    nor g1554(n1430 ,n581 ,n1022);
    nor g1555(n1429 ,n611 ,n1022);
    nor g1556(n1428 ,n596 ,n1022);
    nor g1557(n1427 ,n377 ,n1022);
    nor g1558(n1426 ,n360 ,n1022);
    nor g1559(n1425 ,n561 ,n1022);
    nor g1560(n1424 ,n607 ,n1022);
    nor g1561(n1423 ,n644 ,n1026);
    nor g1562(n1422 ,n402 ,n1026);
    nor g1563(n1421 ,n616 ,n1026);
    nor g1564(n1420 ,n567 ,n1026);
    nor g1565(n1419 ,n681 ,n1026);
    nor g1566(n1418 ,n586 ,n1026);
    nor g1567(n1417 ,n662 ,n1026);
    nor g1568(n1416 ,n695 ,n1026);
    nor g1569(n1415 ,n633 ,n1030);
    nor g1570(n1414 ,n370 ,n1012);
    nor g1571(n1413 ,n613 ,n1030);
    nor g1572(n1412 ,n371 ,n1030);
    nor g1573(n1411 ,n601 ,n1028);
    nor g1574(n1410 ,n392 ,n1030);
    nor g1575(n1409 ,n677 ,n1030);
    nor g1576(n1408 ,n374 ,n1030);
    nor g1577(n1407 ,n658 ,n1024);
    nor g1578(n1406 ,n338 ,n1016);
    nor g1579(n1405 ,n404 ,n1016);
    nor g1580(n1404 ,n623 ,n1016);
    nor g1581(n1403 ,n326 ,n1016);
    nor g1582(n1402 ,n336 ,n1016);
    nor g1583(n1401 ,n669 ,n1016);
    nor g1584(n1400 ,n411 ,n1016);
    nor g1585(n1399 ,n583 ,n1032);
    nor g1586(n1398 ,n368 ,n1032);
    nor g1587(n1397 ,n673 ,n1032);
    nor g1588(n1396 ,n688 ,n1032);
    nor g1589(n1395 ,n617 ,n1032);
    nor g1590(n1394 ,n322 ,n1032);
    nor g1591(n1393 ,n417 ,n1032);
    nor g1592(n1392 ,n614 ,n1032);
    nor g1593(n1391 ,n541 ,n1034);
    nor g1594(n1390 ,n637 ,n1012);
    nor g1595(n1389 ,n651 ,n1034);
    nor g1596(n1388 ,n430 ,n1034);
    nor g1597(n1387 ,n577 ,n1034);
    nor g1598(n1386 ,n652 ,n1034);
    nor g1599(n1385 ,n570 ,n1006);
    nor g1600(n1384 ,n343 ,n1006);
    nor g1601(n1383 ,n436 ,n1006);
    nor g1602(n1382 ,n363 ,n1006);
    nor g1603(n1381 ,n388 ,n1006);
    nor g1604(n1380 ,n397 ,n1006);
    nor g1605(n1379 ,n592 ,n1018);
    nor g1606(n1378 ,n544 ,n1018);
    nor g1607(n1377 ,n612 ,n1018);
    nor g1608(n1376 ,n547 ,n1024);
    nor g1609(n1375 ,n345 ,n1018);
    nor g1610(n1374 ,n622 ,n1018);
    nor g1611(n1373 ,n394 ,n1018);
    nor g1612(n1372 ,n619 ,n1018);
    nor g1613(n1371 ,n597 ,n1008);
    nor g1614(n1370 ,n552 ,n1008);
    nor g1615(n1369 ,n572 ,n1008);
    nor g1616(n1368 ,n571 ,n1008);
    nor g1617(n1367 ,n419 ,n1008);
    nor g1618(n1366 ,n340 ,n1008);
    nor g1619(n1365 ,n600 ,n1024);
    nor g1620(n1364 ,n691 ,n1024);
    nor g1621(n1363 ,n564 ,n1024);
    nor g1622(n1362 ,n414 ,n1024);
    nor g1623(n1361 ,n373 ,n1024);
    nor g1624(n1360 ,n625 ,n1024);
    nor g1625(n1359 ,n557 ,n1014);
    nor g1626(n1358 ,n539 ,n1028);
    nor g1627(n1357 ,n429 ,n1028);
    nor g1628(n1356 ,n587 ,n1028);
    nor g1629(n1355 ,n425 ,n1028);
    nor g1630(n1354 ,n341 ,n1028);
    nor g1631(n1353 ,n685 ,n1028);
    nor g1632(n1352 ,n648 ,n1014);
    nor g1633(n1351 ,n405 ,n1014);
    nor g1634(n1350 ,n659 ,n1014);
    nor g1635(n1349 ,n508 ,n1039);
    nor g1636(n1348 ,n509 ,n1039);
    nor g1637(n1347 ,n304 ,n1038);
    nor g1638(n1346 ,n292 ,n1011);
    or g1639(n1345 ,n770 ,n946);
    nor g1640(n1344 ,n299 ,n1047);
    nor g1641(n1343 ,n296 ,n1013);
    nor g1642(n1342 ,n298 ,n1013);
    nor g1643(n1341 ,n295 ,n1019);
    nor g1644(n1340 ,n297 ,n1019);
    nor g1645(n1339 ,n293 ,n1019);
    nor g1646(n1338 ,n294 ,n1019);
    nor g1647(n1337 ,n296 ,n1019);
    nor g1648(n1336 ,n298 ,n1019);
    nor g1649(n1335 ,n295 ,n1011);
    nor g1650(n1334 ,n293 ,n1011);
    or g1651(n1516 ,n515 ,n1036);
    or g1652(n1515 ,n705 ,n948);
    not g1653(n1333 ,n1332);
    not g1654(n1331 ,n1330);
    not g1655(n1322 ,n1323);
    xnor g1656(n1321 ,n928 ,n59[0]);
    nor g1657(n1320 ,n296 ,n1011);
    nor g1658(n1319 ,n297 ,n1033);
    nor g1659(n1318 ,n294 ,n1011);
    nor g1660(n1317 ,n295 ,n1021);
    nor g1661(n1316 ,n291 ,n1021);
    nor g1662(n1315 ,n297 ,n1021);
    nor g1663(n1314 ,n293 ,n1021);
    nor g1664(n1313 ,n291 ,n1015);
    nor g1665(n1312 ,n294 ,n1021);
    nor g1666(n1311 ,n292 ,n1021);
    nor g1667(n1310 ,n296 ,n1021);
    nor g1668(n1309 ,n298 ,n1021);
    nor g1669(n1308 ,n295 ,n1025);
    nor g1670(n1307 ,n291 ,n1025);
    nor g1671(n1306 ,n297 ,n1011);
    nor g1672(n1305 ,n298 ,n1005);
    nor g1673(n1304 ,n297 ,n1025);
    nor g1674(n1303 ,n293 ,n1025);
    nor g1675(n1302 ,n294 ,n1025);
    nor g1676(n1301 ,n292 ,n1025);
    nor g1677(n1300 ,n296 ,n1025);
    nor g1678(n1299 ,n298 ,n1025);
    nor g1679(n1298 ,n295 ,n1029);
    nor g1680(n1297 ,n291 ,n1029);
    nor g1681(n1296 ,n297 ,n1029);
    nor g1682(n1295 ,n293 ,n1029);
    nor g1683(n1294 ,n294 ,n1029);
    nor g1684(n1293 ,n292 ,n1029);
    nor g1685(n1292 ,n296 ,n1029);
    nor g1686(n1291 ,n298 ,n1029);
    nor g1687(n1290 ,n295 ,n1015);
    nor g1688(n1289 ,n297 ,n1015);
    nor g1689(n1288 ,n293 ,n1015);
    nor g1690(n1287 ,n294 ,n1015);
    nor g1691(n1286 ,n292 ,n1015);
    nor g1692(n1285 ,n296 ,n1015);
    nor g1693(n1284 ,n291 ,n1011);
    nor g1694(n1283 ,n298 ,n1015);
    nor g1695(n1282 ,n295 ,n1031);
    nor g1696(n1281 ,n291 ,n1031);
    nor g1697(n1280 ,n297 ,n1031);
    nor g1698(n1279 ,n293 ,n1031);
    nor g1699(n1278 ,n294 ,n1031);
    nor g1700(n1277 ,n292 ,n1031);
    nor g1701(n1276 ,n296 ,n1031);
    nor g1702(n1275 ,n298 ,n1031);
    nor g1703(n1274 ,n295 ,n1033);
    nor g1704(n1273 ,n291 ,n1033);
    nor g1705(n1272 ,n293 ,n1033);
    nor g1706(n1271 ,n294 ,n1033);
    nor g1707(n1270 ,n292 ,n1033);
    nor g1708(n1269 ,n296 ,n1033);
    nor g1709(n1268 ,n298 ,n1033);
    nor g1710(n1267 ,n295 ,n1005);
    nor g1711(n1266 ,n291 ,n1005);
    nor g1712(n1265 ,n297 ,n1005);
    nor g1713(n1264 ,n293 ,n1005);
    nor g1714(n1263 ,n294 ,n1005);
    nor g1715(n1262 ,n292 ,n1005);
    nor g1716(n1261 ,n296 ,n1005);
    nor g1717(n1260 ,n295 ,n1017);
    nor g1718(n1259 ,n291 ,n1017);
    nor g1719(n1258 ,n297 ,n1017);
    nor g1720(n1257 ,n293 ,n1017);
    nor g1721(n1256 ,n294 ,n1017);
    nor g1722(n1255 ,n292 ,n1017);
    nor g1723(n1254 ,n296 ,n1017);
    nor g1724(n1253 ,n298 ,n1017);
    nor g1725(n1252 ,n292 ,n1019);
    nor g1726(n1251 ,n295 ,n1007);
    nor g1727(n1250 ,n291 ,n1007);
    nor g1728(n1249 ,n297 ,n1007);
    nor g1729(n1248 ,n293 ,n1007);
    nor g1730(n1247 ,n294 ,n1007);
    nor g1731(n1246 ,n292 ,n1007);
    nor g1732(n1245 ,n296 ,n1007);
    nor g1733(n1244 ,n298 ,n1007);
    nor g1734(n1243 ,n295 ,n1023);
    nor g1735(n1242 ,n291 ,n1023);
    nor g1736(n1241 ,n297 ,n1023);
    nor g1737(n1240 ,n293 ,n1023);
    nor g1738(n1239 ,n294 ,n1023);
    nor g1739(n1238 ,n292 ,n1023);
    nor g1740(n1237 ,n296 ,n1023);
    nor g1741(n1236 ,n298 ,n1023);
    nor g1742(n1235 ,n295 ,n1027);
    nor g1743(n1234 ,n291 ,n1027);
    nor g1744(n1233 ,n297 ,n1027);
    nor g1745(n1232 ,n293 ,n1027);
    nor g1746(n1231 ,n294 ,n1027);
    nor g1747(n1230 ,n292 ,n1027);
    nor g1748(n1229 ,n296 ,n1027);
    nor g1749(n1228 ,n298 ,n1027);
    nor g1750(n1227 ,n295 ,n1013);
    nor g1751(n1226 ,n291 ,n1013);
    nor g1752(n1225 ,n297 ,n1013);
    nor g1753(n1224 ,n293 ,n1013);
    nor g1754(n1223 ,n294 ,n1013);
    nor g1755(n1222 ,n292 ,n1013);
    nor g1756(n1221 ,n296 ,n1003);
    nor g1757(n1220 ,n294 ,n1003);
    nor g1758(n1219 ,n295 ,n1003);
    nor g1759(n1218 ,n291 ,n1003);
    nor g1760(n1217 ,n293 ,n1003);
    nor g1761(n1216 ,n292 ,n1003);
    nor g1762(n1215 ,n298 ,n1003);
    nor g1763(n1214 ,n297 ,n1003);
    nor g1764(n1213 ,n293 ,n1009);
    nor g1765(n1212 ,n499 ,n947);
    nor g1766(n1211 ,n725 ,n1037);
    or g1767(n1210 ,n968 ,n970);
    nor g1768(n1209 ,n791 ,n944);
    or g1769(n1208 ,n987 ,n1100);
    or g1770(n1207 ,n974 ,n1075);
    or g1771(n1206 ,n1108 ,n998);
    or g1772(n1205 ,n1096 ,n1122);
    or g1773(n1204 ,n1090 ,n1128);
    or g1774(n1203 ,n1088 ,n1135);
    or g1775(n1202 ,n1134 ,n1136);
    or g1776(n1201 ,n1094 ,n978);
    or g1777(n1200 ,n1099 ,n972);
    or g1778(n1199 ,n975 ,n1114);
    or g1779(n1198 ,n986 ,n985);
    or g1780(n1197 ,n1061 ,n1124);
    or g1781(n1196 ,n1121 ,n967);
    or g1782(n1195 ,n1087 ,n1093);
    nor g1783(n1194 ,n710 ,n945);
    or g1784(n1193 ,n1097 ,n1104);
    or g1785(n1192 ,n1086 ,n1111);
    or g1786(n1191 ,n1110 ,n1076);
    or g1787(n1190 ,n1138 ,n1127);
    or g1788(n1189 ,n992 ,n1089);
    or g1789(n1188 ,n1084 ,n1060);
    or g1790(n1187 ,n981 ,n1137);
    or g1791(n1186 ,n17[0] ,n1045);
    or g1792(n1185 ,n1113 ,n1120);
    or g1793(n1184 ,n973 ,n1118);
    or g1794(n1183 ,n1126 ,n1119);
    or g1795(n1182 ,n1092 ,n1058);
    or g1796(n1181 ,n1139 ,n1106);
    or g1797(n1180 ,n1109 ,n1117);
    or g1798(n1179 ,n971 ,n989);
    or g1799(n1178 ,n1103 ,n1130);
    or g1800(n1177 ,n1116 ,n1102);
    or g1801(n1176 ,n977 ,n1085);
    or g1802(n1175 ,n1083 ,n1082);
    or g1803(n1174 ,n1081 ,n1080);
    or g1804(n1173 ,n1079 ,n1077);
    or g1805(n1172 ,n980 ,n1073);
    or g1806(n1171 ,n1074 ,n1072);
    or g1807(n1170 ,n1071 ,n1066);
    or g1808(n1169 ,n1070 ,n1069);
    or g1809(n1168 ,n1068 ,n1067);
    or g1810(n1167 ,n1065 ,n1064);
    or g1811(n1166 ,n1054 ,n1063);
    or g1812(n1165 ,n1059 ,n1057);
    or g1813(n1164 ,n1056 ,n1055);
    or g1814(n1163 ,n1052 ,n1131);
    nor g1815(n1162 ,n906 ,n943);
    or g1816(n1161 ,n1053 ,n1051);
    nor g1817(n1160 ,n905 ,n957);
    nor g1818(n1159 ,n902 ,n956);
    nor g1819(n1158 ,n909 ,n950);
    or g1820(n1157 ,n994 ,n1050);
    nor g1821(n1156 ,n904 ,n955);
    or g1822(n1155 ,n1049 ,n1095);
    nor g1823(n1154 ,n903 ,n1002);
    nor g1824(n1153 ,n901 ,n953);
    nor g1825(n1152 ,n900 ,n952);
    or g1826(n1151 ,n954 ,n1001);
    nor g1827(n1150 ,n908 ,n951);
    or g1828(n1149 ,n996 ,n999);
    nor g1829(n1148 ,n910 ,n958);
    or g1830(n1147 ,n1000 ,n997);
    nor g1831(n1146 ,n899 ,n949);
    or g1832(n1145 ,n995 ,n991);
    or g1833(n1144 ,n976 ,n1107);
    or g1834(n1143 ,n990 ,n988);
    nor g1835(n1142 ,n62[2] ,n1043);
    or g1836(n1141 ,n993 ,n1123);
    or g1837(n1140 ,n982 ,n983);
    nor g1838(n1332 ,n826 ,n932);
    nor g1839(n1330 ,n793 ,n1040);
    or g1840(n1329 ,n59[3] ,n1036);
    or g1841(n1328 ,n278 ,n1041);
    or g1842(n1327 ,n279 ,n934);
    or g1843(n1325 ,n279 ,n1040);
    or g1844(n1324 ,n921 ,n1039);
    nor g1845(n1323 ,n2653 ,n1040);
    nor g1846(n1139 ,n660 ,n916);
    nor g1847(n1138 ,n361 ,n926);
    nor g1848(n1137 ,n383 ,n917);
    nor g1849(n1136 ,n663 ,n919);
    nor g1850(n1135 ,n609 ,n883);
    nor g1851(n1134 ,n410 ,n920);
    nor g1852(n1133 ,n424 ,n922);
    nor g1853(n1132 ,n380 ,n924);
    nor g1854(n1131 ,n582 ,n883);
    nor g1855(n1130 ,n670 ,n919);
    nor g1856(n1129 ,n655 ,n924);
    nor g1857(n1128 ,n690 ,n917);
    nor g1858(n1127 ,n426 ,n888);
    nor g1859(n1126 ,n324 ,n925);
    nor g1860(n1125 ,n428 ,n924);
    nor g1861(n1124 ,n335 ,n919);
    nor g1862(n1123 ,n439 ,n883);
    nor g1863(n1122 ,n578 ,n917);
    nor g1864(n1121 ,n537 ,n916);
    nor g1865(n1120 ,n418 ,n885);
    nor g1866(n1119 ,n339 ,n883);
    nor g1867(n1118 ,n560 ,n883);
    nor g1868(n1117 ,n696 ,n885);
    nor g1869(n1116 ,n684 ,n926);
    nor g1870(n1115 ,n573 ,n922);
    nor g1871(n1114 ,n589 ,n888);
    nor g1872(n1113 ,n364 ,n884);
    nor g1873(n1112 ,n441 ,n924);
    nor g1874(n1111 ,n337 ,n886);
    nor g1875(n1110 ,n349 ,n887);
    nor g1876(n1109 ,n386 ,n884);
    nor g1877(n1108 ,n412 ,n926);
    nor g1878(n1107 ,n344 ,n886);
    nor g1879(n1106 ,n689 ,n923);
    nor g1880(n1105 ,n545 ,n922);
    nor g1881(n1104 ,n640 ,n923);
    nor g1882(n1103 ,n346 ,n920);
    nor g1883(n1102 ,n382 ,n888);
    nor g1884(n1101 ,n331 ,n924);
    nor g1885(n1100 ,n548 ,n886);
    nor g1886(n1099 ,n591 ,n887);
    nor g1887(n1098 ,n590 ,n922);
    nor g1888(n1097 ,n378 ,n916);
    nor g1889(n1096 ,n643 ,n918);
    nor g1890(n1095 ,n683 ,n888);
    nor g1891(n1094 ,n372 ,n926);
    nor g1892(n1093 ,n615 ,n917);
    nor g1893(n1092 ,n551 ,n884);
    nor g1894(n1091 ,n549 ,n922);
    nor g1895(n1090 ,n671 ,n918);
    nor g1896(n1089 ,n389 ,n885);
    nor g1897(n1088 ,n396 ,n925);
    nor g1898(n1087 ,n393 ,n918);
    nor g1899(n1086 ,n442 ,n887);
    nor g1900(n1085 ,n351 ,n917);
    nor g1901(n1084 ,n438 ,n884);
    nor g1902(n1083 ,n321 ,n920);
    nor g1903(n1082 ,n327 ,n919);
    nor g1904(n1081 ,n536 ,n918);
    nor g1905(n1080 ,n558 ,n917);
    nor g1906(n1079 ,n427 ,n925);
    nor g1907(n1078 ,n603 ,n922);
    nor g1908(n1077 ,n585 ,n883);
    nor g1909(n1076 ,n606 ,n886);
    nor g1910(n1075 ,n657 ,n919);
    nor g1911(n1074 ,n647 ,n916);
    nor g1912(n1073 ,n635 ,n923);
    nor g1913(n1072 ,n568 ,n923);
    nor g1914(n1071 ,n329 ,n920);
    nor g1915(n1070 ,n668 ,n926);
    nor g1916(n1069 ,n674 ,n888);
    nor g1917(n1068 ,n649 ,n887);
    nor g1918(n1067 ,n636 ,n886);
    nor g1919(n1066 ,n406 ,n919);
    nor g1920(n1065 ,n367 ,n884);
    nor g1921(n1064 ,n432 ,n885);
    nor g1922(n1063 ,n628 ,n917);
    nor g1923(n1062 ,n574 ,n924);
    nor g1924(n1061 ,n415 ,n920);
    nor g1925(n1060 ,n422 ,n885);
    nor g1926(n1059 ,n318 ,n920);
    nor g1927(n1058 ,n348 ,n885);
    nor g1928(n1057 ,n362 ,n919);
    nor g1929(n1056 ,n630 ,n918);
    nor g1930(n1055 ,n580 ,n917);
    nor g1931(n1054 ,n385 ,n918);
    nor g1932(n1053 ,n694 ,n925);
    nor g1933(n1052 ,n624 ,n925);
    nor g1934(n1051 ,n653 ,n883);
    nor g1935(n1050 ,n593 ,n923);
    nor g1936(n1049 ,n403 ,n926);
    not g1937(n1048 ,n1047);
    not g1938(n1046 ,n1045);
    not g1939(n1044 ,n1043);
    not g1940(n1041 ,n1040);
    not g1941(n1038 ,n1037);
    not g1942(n1033 ,n1034);
    not g1943(n1031 ,n1032);
    not g1944(n1029 ,n1030);
    not g1945(n1027 ,n1028);
    not g1946(n1025 ,n1026);
    not g1947(n1023 ,n1024);
    not g1948(n1021 ,n1022);
    not g1949(n1019 ,n1020);
    not g1950(n1017 ,n1018);
    not g1951(n1015 ,n1016);
    not g1952(n1013 ,n1014);
    not g1953(n1011 ,n1012);
    not g1954(n1009 ,n1010);
    not g1955(n1007 ,n1008);
    not g1956(n1005 ,n1006);
    not g1957(n1003 ,n1004);
    nor g1958(n1002 ,n482 ,n882);
    nor g1959(n1001 ,n350 ,n886);
    nor g1960(n1000 ,n384 ,n884);
    nor g1961(n999 ,n697 ,n923);
    nor g1962(n998 ,n631 ,n888);
    nor g1963(n997 ,n692 ,n885);
    nor g1964(n996 ,n400 ,n916);
    nor g1965(n995 ,n413 ,n926);
    nor g1966(n994 ,n654 ,n916);
    nor g1967(n993 ,n665 ,n925);
    nor g1968(n992 ,n576 ,n884);
    nor g1969(n991 ,n559 ,n888);
    nor g1970(n990 ,n584 ,n887);
    nor g1971(n989 ,n579 ,n883);
    nor g1972(n988 ,n682 ,n886);
    nor g1973(n987 ,n398 ,n887);
    nor g1974(n986 ,n645 ,n884);
    nor g1975(n985 ,n599 ,n885);
    nor g1976(n984 ,n538 ,n924);
    nor g1977(n983 ,n605 ,n919);
    nor g1978(n982 ,n409 ,n920);
    nor g1979(n981 ,n358 ,n918);
    nor g1980(n980 ,n627 ,n916);
    nor g1981(n979 ,n352 ,n924);
    nor g1982(n978 ,n650 ,n888);
    nor g1983(n977 ,n408 ,n918);
    nor g1984(n976 ,n354 ,n887);
    nor g1985(n975 ,n676 ,n926);
    nor g1986(n974 ,n319 ,n920);
    nor g1987(n973 ,n540 ,n925);
    nor g1988(n972 ,n440 ,n886);
    nor g1989(n971 ,n334 ,n925);
    nor g1990(n970 ,n332 ,n923);
    nor g1991(n969 ,n604 ,n922);
    nor g1992(n968 ,n687 ,n916);
    nor g1993(n967 ,n608 ,n923);
    nor g1994(n966 ,n433 ,n915);
    nor g1995(n965 ,n434 ,n915);
    nor g1996(n964 ,n379 ,n915);
    nor g1997(n963 ,n399 ,n915);
    nor g1998(n962 ,n562 ,n915);
    nor g1999(n961 ,n641 ,n915);
    nor g2000(n960 ,n357 ,n915);
    nor g2001(n959 ,n375 ,n915);
    nor g2002(n958 ,n491 ,n882);
    nor g2003(n957 ,n452 ,n882);
    nor g2004(n956 ,n479 ,n882);
    nor g2005(n955 ,n488 ,n882);
    nor g2006(n954 ,n661 ,n887);
    nor g2007(n953 ,n446 ,n882);
    nor g2008(n952 ,n464 ,n882);
    nor g2009(n951 ,n480 ,n882);
    nor g2010(n950 ,n489 ,n882);
    nor g2011(n949 ,n459 ,n882);
    or g2012(n948 ,n879 ,n896);
    nor g2013(n947 ,n17[2] ,n907);
    or g2014(n946 ,n856 ,n912);
    nor g2015(n945 ,n62[2] ,n911);
    or g2016(n944 ,n17[1] ,n870);
    nor g2017(n943 ,n40[0] ,n882);
    nor g2018(n942 ,n286 ,n866);
    nor g2019(n941 ,n283 ,n874);
    nor g2020(n940 ,n284 ,n867);
    nor g2021(n939 ,n280 ,n876);
    nor g2022(n938 ,n284 ,n864);
    nor g2023(n937 ,n285 ,n869);
    nor g2024(n936 ,n285 ,n865);
    nor g2025(n935 ,n281 ,n873);
    nor g2026(n934 ,n897 ,n896);
    nor g2027(n933 ,n878 ,n877);
    nor g2028(n932 ,n844 ,n868);
    nor g2029(n1047 ,n784 ,n895);
    nor g2030(n1045 ,n930 ,n875);
    nor g2031(n1043 ,n928 ,n895);
    or g2032(n1042 ,n747 ,n914);
    nor g2033(n1040 ,n19[4] ,n931);
    or g2034(n1039 ,n279 ,n928);
    nor g2035(n1037 ,n783 ,n928);
    or g2036(n1036 ,n286 ,n927);
    or g2037(n1035 ,n286 ,n893);
    nor g2038(n1034 ,n720 ,n889);
    nor g2039(n1032 ,n720 ,n890);
    nor g2040(n1030 ,n712 ,n890);
    nor g2041(n1028 ,n712 ,n891);
    nor g2042(n1026 ,n714 ,n889);
    nor g2043(n1024 ,n714 ,n929);
    nor g2044(n1022 ,n714 ,n890);
    nor g2045(n1020 ,n720 ,n891);
    nor g2046(n1018 ,n750 ,n889);
    nor g2047(n1016 ,n712 ,n889);
    nor g2048(n1014 ,n712 ,n929);
    nor g2049(n1012 ,n720 ,n929);
    nor g2050(n1010 ,n750 ,n891);
    nor g2051(n1008 ,n714 ,n891);
    nor g2052(n1006 ,n750 ,n890);
    nor g2053(n1004 ,n750 ,n929);
    not g2054(n931 ,n930);
    not g2055(n927 ,n928);
    not g2056(n922 ,n921);
    not g2057(n915 ,n914);
    nor g2058(n913 ,n304 ,n861);
    nor g2059(n912 ,n543 ,n863);
    nor g2060(n911 ,n300 ,n838);
    nor g2061(n910 ,n518 ,n829);
    nor g2062(n909 ,n526 ,n829);
    nor g2063(n908 ,n521 ,n829);
    nor g2064(n907 ,n313 ,n817);
    nor g2065(n906 ,n311 ,n829);
    nor g2066(n905 ,n531 ,n829);
    nor g2067(n904 ,n520 ,n829);
    nor g2068(n903 ,n535 ,n829);
    nor g2069(n902 ,n312 ,n829);
    nor g2070(n901 ,n314 ,n829);
    nor g2071(n900 ,n315 ,n829);
    nor g2072(n899 ,n516 ,n829);
    nor g2073(n898 ,n511 ,n862);
    or g2074(n897 ,n300 ,n827);
    nor g2075(n930 ,n498 ,n809);
    or g2076(n929 ,n301 ,n860);
    nor g2077(n928 ,n2597 ,n813);
    or g2078(n926 ,n722 ,n859);
    or g2079(n925 ,n718 ,n858);
    or g2080(n924 ,n722 ,n831);
    or g2081(n923 ,n711 ,n831);
    nor g2082(n921 ,n300 ,n863);
    or g2083(n920 ,n751 ,n831);
    or g2084(n919 ,n711 ,n858);
    or g2085(n918 ,n751 ,n859);
    or g2086(n917 ,n718 ,n831);
    or g2087(n916 ,n718 ,n859);
    nor g2088(n914 ,n751 ,n858);
    not g2089(n894 ,n893);
    or g2090(n880 ,n843 ,n836);
    nor g2091(n879 ,n62[2] ,n838);
    or g2092(n878 ,n17[1] ,n811);
    nor g2093(n877 ,n17[2] ,n834);
    nor g2094(n876 ,n821 ,n850);
    nor g2095(n875 ,n728 ,n812);
    nor g2096(n874 ,n822 ,n851);
    nor g2097(n873 ,n824 ,n839);
    nor g2098(n872 ,n19[4] ,n862);
    nor g2099(n871 ,n58[4] ,n861);
    nor g2100(n870 ,n17[2] ,n835);
    nor g2101(n869 ,n823 ,n841);
    or g2102(n868 ,n17[1] ,n832);
    nor g2103(n867 ,n818 ,n846);
    nor g2104(n866 ,n820 ,n840);
    nor g2105(n865 ,n825 ,n814);
    nor g2106(n864 ,n819 ,n847);
    nor g2107(n896 ,n299 ,n810);
    nor g2108(n895 ,n772 ,n849);
    nor g2109(n893 ,n699 ,n816);
    nor g2110(n892 ,n17[1] ,n833);
    or g2111(n891 ,n60[0] ,n860);
    or g2112(n890 ,n60[3] ,n837);
    or g2113(n889 ,n60[3] ,n842);
    or g2114(n888 ,n711 ,n859);
    or g2115(n887 ,n751 ,n830);
    or g2116(n886 ,n718 ,n830);
    or g2117(n885 ,n711 ,n830);
    or g2118(n884 ,n722 ,n830);
    or g2119(n883 ,n722 ,n858);
    or g2120(n882 ,n2655 ,n828);
    nor g2121(n857 ,n507 ,n783);
    nor g2122(n856 ,n672 ,n787);
    nor g2123(n855 ,n468 ,n782);
    nor g2124(n854 ,n449 ,n782);
    nor g2125(n853 ,n476 ,n782);
    nor g2126(n852 ,n457 ,n782);
    nor g2127(n851 ,n494 ,n780);
    nor g2128(n850 ,n288 ,n780);
    or g2129(n849 ,n300 ,n796);
    nor g2130(n848 ,n306 ,n783);
    nor g2131(n847 ,n290 ,n780);
    nor g2132(n846 ,n305 ,n780);
    nor g2133(n845 ,n503 ,n783);
    nor g2134(n844 ,n328 ,n792);
    nor g2135(n843 ,n301 ,n783);
    or g2136(n842 ,n301 ,n782);
    nor g2137(n841 ,n496 ,n780);
    nor g2138(n840 ,n495 ,n780);
    nor g2139(n839 ,n289 ,n780);
    or g2140(n863 ,n278 ,n779);
    or g2141(n862 ,n704 ,n769);
    or g2142(n861 ,n702 ,n766);
    or g2143(n860 ,n306 ,n782);
    or g2144(n859 ,n303 ,n797);
    or g2145(n858 ,n303 ,n808);
    not g2146(n837 ,n836);
    not g2147(n835 ,n834);
    not g2148(n833 ,n832);
    not g2149(n829 ,n828);
    nor g2150(n827 ,n755 ,n778);
    nor g2151(n826 ,n499 ,n763);
    nor g2152(n825 ,n497 ,n781);
    nor g2153(n824 ,n496 ,n781);
    nor g2154(n823 ,n287 ,n781);
    nor g2155(n822 ,n290 ,n781);
    nor g2156(n821 ,n494 ,n781);
    nor g2157(n820 ,n288 ,n781);
    nor g2158(n819 ,n289 ,n781);
    nor g2159(n818 ,n495 ,n781);
    nor g2160(n817 ,n17[0] ,n807);
    nor g2161(n816 ,n774 ,n773);
    or g2162(n815 ,n764 ,n775);
    nor g2163(n814 ,n287 ,n780);
    or g2164(n813 ,n4 ,n785);
    or g2165(n812 ,n698 ,n788);
    nor g2166(n811 ,n727 ,n789);
    nor g2167(n810 ,n709 ,n795);
    or g2168(n809 ,n17[1] ,n790);
    nor g2169(n838 ,n724 ,n804);
    nor g2170(n836 ,n60[0] ,n782);
    nor g2171(n834 ,n771 ,n788);
    nor g2172(n832 ,n2 ,n768);
    or g2173(n831 ,n37[2] ,n808);
    or g2174(n830 ,n37[2] ,n797);
    or g2175(n828 ,n786 ,n784);
    nor g2176(n806 ,n420 ,n708);
    nor g2177(n805 ,n390 ,n708);
    nor g2178(n804 ,n310 ,n745);
    nor g2179(n803 ,n678 ,n708);
    nor g2180(n802 ,n675 ,n708);
    nor g2181(n801 ,n639 ,n708);
    nor g2182(n800 ,n330 ,n708);
    nor g2183(n799 ,n309 ,n708);
    nor g2184(n798 ,n376 ,n708);
    or g2185(n808 ,n309 ,n747);
    nor g2186(n807 ,n523 ,n746);
    not g2187(n796 ,n795);
    not g2188(n794 ,n793);
    not g2189(n792 ,n791);
    not g2190(n790 ,n789);
    not g2191(n787 ,n786);
    not g2192(n785 ,n784);
    not g2193(n780 ,n781);
    or g2194(n779 ,n62[2] ,n724);
    or g2195(n778 ,n62[2] ,n723);
    nor g2196(n777 ,n303 ,n708);
    nor g2197(n776 ,n302 ,n708);
    nor g2198(n775 ,n502 ,n708);
    nor g2199(n774 ,n17[2] ,n706);
    or g2200(n773 ,n17[1] ,n726);
    or g2201(n772 ,n299 ,n709);
    nor g2202(n771 ,n500 ,n753);
    or g2203(n770 ,n278 ,n710);
    or g2204(n769 ,n278 ,n703);
    or g2205(n768 ,n17[2] ,n754);
    nor g2206(n767 ,n499 ,n760);
    or g2207(n766 ,n58[1] ,n725);
    nor g2208(n765 ,n626 ,n708);
    nor g2209(n764 ,n37[0] ,n747);
    nor g2210(n763 ,n17[0] ,n761);
    or g2211(n762 ,n62[2] ,n756);
    or g2212(n797 ,n37[3] ,n747);
    nor g2213(n795 ,n41[1] ,n701);
    nor g2214(n793 ,n17[0] ,n728);
    nor g2215(n791 ,n498 ,n752);
    nor g2216(n789 ,n2646 ,n752);
    nor g2217(n788 ,n305 ,n753);
    nor g2218(n786 ,n299 ,n710);
    nor g2219(n784 ,n62[2] ,n709);
    or g2220(n783 ,n278 ,n757);
    or g2221(n782 ,n278 ,n758);
    nor g2222(n781 ,n752 ,n729);
    not g2223(n761 ,n760);
    not g2224(n758 ,n757);
    not g2225(n756 ,n755);
    not g2226(n754 ,n753);
    or g2227(n746 ,n512 ,n317);
    or g2228(n745 ,n510 ,n514);
    nor g2229(n744 ,n517 ,n283);
    nor g2230(n743 ,n311 ,n284);
    nor g2231(n742 ,n520 ,n280);
    nor g2232(n741 ,n524 ,n281);
    nor g2233(n740 ,n312 ,n284);
    nor g2234(n739 ,n518 ,n283);
    nor g2235(n738 ,n314 ,n285);
    nor g2236(n737 ,n526 ,n282);
    nor g2237(n736 ,n530 ,n283);
    nor g2238(n735 ,n315 ,n282);
    nor g2239(n734 ,n516 ,n283);
    nor g2240(n733 ,n521 ,n281);
    nor g2241(n732 ,n535 ,n280);
    nor g2242(n731 ,n531 ,n281);
    nor g2243(n730 ,n533 ,n282);
    nor g2244(n760 ,n313 ,n17[2]);
    nor g2245(n759 ,n575 ,n282);
    nor g2246(n757 ,n320 ,n58[4]);
    nor g2247(n755 ,n308 ,n62[1]);
    nor g2248(n753 ,n500 ,n2596);
    or g2249(n752 ,n313 ,n17[0]);
    or g2250(n751 ,n502 ,n302);
    or g2251(n750 ,n507 ,n503);
    or g2252(n749 ,n508 ,n509);
    or g2253(n748 ,n504 ,n506);
    or g2254(n747 ,n279 ,n316);
    not g2255(n727 ,n726);
    not g2256(n724 ,n723);
    not g2257(n709 ,n710);
    or g2258(n707 ,n307 ,n62[2]);
    nor g2259(n706 ,n305 ,n17[0]);
    or g2260(n705 ,n279 ,n300);
    or g2261(n704 ,n19[2] ,n19[3]);
    or g2262(n703 ,n19[0] ,n19[1]);
    or g2263(n702 ,n58[2] ,n58[3]);
    or g2264(n701 ,n41[0] ,n41[2]);
    or g2265(n700 ,n278 ,n2652);
    nor g2266(n699 ,n499 ,n498);
    nor g2267(n698 ,n500 ,n2);
    or g2268(n729 ,n499 ,n17[2]);
    or g2269(n728 ,n17[1] ,n17[2]);
    nor g2270(n726 ,n498 ,n17[0]);
    or g2271(n725 ,n279 ,n58[0]);
    nor g2272(n723 ,n307 ,n62[0]);
    or g2273(n722 ,n502 ,n37[1]);
    or g2274(n721 ,n508 ,n59[2]);
    or g2275(n720 ,n503 ,n60[1]);
    or g2276(n719 ,n59[1] ,n59[2]);
    or g2277(n718 ,n302 ,n37[0]);
    or g2278(n717 ,n38[1] ,n38[2]);
    or g2279(n716 ,n509 ,n59[1]);
    or g2280(n715 ,n506 ,n38[1]);
    or g2281(n714 ,n60[1] ,n60[2]);
    or g2282(n713 ,n504 ,n38[2]);
    or g2283(n712 ,n507 ,n60[2]);
    or g2284(n711 ,n37[0] ,n37[1]);
    nor g2285(n710 ,n62[0] ,n62[1]);
    or g2286(n708 ,n279 ,n2653);
    not g2287(n697 ,n29[0]);
    not g2288(n696 ,n21[1]);
    not g2289(n695 ,n43[7]);
    not g2290(n694 ,n35[7]);
    not g2291(n693 ,n54[2]);
    not g2292(n692 ,n21[7]);
    not g2293(n691 ,n51[1]);
    not g2294(n690 ,n31[3]);
    not g2295(n689 ,n29[3]);
    not g2296(n688 ,n46[3]);
    not g2297(n687 ,n27[2]);
    not g2298(n686 ,n20[5]);
    not g2299(n685 ,n52[7]);
    not g2300(n684 ,n26[4]);
    not g2301(n683 ,n25[7]);
    not g2302(n682 ,n23[0]);
    not g2303(n681 ,n43[4]);
    not g2304(n680 ,n56[3]);
    not g2305(n679 ,n53[7]);
    not g2306(n678 ,n12[1]);
    not g2307(n677 ,n44[5]);
    not g2308(n676 ,n26[5]);
    not g2309(n675 ,n12[0]);
    not g2310(n674 ,n25[6]);
    not g2311(n673 ,n46[2]);
    not g2312(n672 ,n6);
    not g2313(n671 ,n28[3]);
    not g2314(n670 ,n33[5]);
    not g2315(n669 ,n45[6]);
    not g2316(n668 ,n26[6]);
    not g2317(n667 ,n44[7]);
    not g2318(n666 ,n54[4]);
    not g2319(n665 ,n35[1]);
    not g2320(n664 ,n55[4]);
    not g2321(n663 ,n33[1]);
    not g2322(n662 ,n43[6]);
    not g2323(n661 ,n24[7]);
    not g2324(n660 ,n27[3]);
    not g2325(n659 ,n53[3]);
    not g2326(n658 ,n51[7]);
    not g2327(n657 ,n33[2]);
    not g2328(n656 ,n20[8]);
    not g2329(n655 ,n30[5]);
    not g2330(n654 ,n27[7]);
    not g2331(n653 ,n34[7]);
    not g2332(n652 ,n47[7]);
    not g2333(n651 ,n47[4]);
    not g2334(n650 ,n25[1]);
    not g2335(n649 ,n24[6]);
    not g2336(n648 ,n53[1]);
    not g2337(n647 ,n27[6]);
    not g2338(n646 ,n54[0]);
    not g2339(n645 ,n22[0]);
    not g2340(n644 ,n43[0]);
    not g2341(n643 ,n28[2]);
    not g2342(n642 ,n20[12]);
    not g2343(n641 ,n36[7]);
    not g2344(n640 ,n29[4]);
    not g2345(n639 ,n12[2]);
    not g2346(n638 ,n20[9]);
    not g2347(n637 ,n55[0]);
    not g2348(n636 ,n23[6]);
    not g2349(n635 ,n29[1]);
    not g2350(n634 ,n49[4]);
    not g2351(n633 ,n44[0]);
    not g2352(n632 ,n53[0]);
    not g2353(n631 ,n25[2]);
    not g2354(n630 ,n28[7]);
    not g2355(n629 ,n20[6]);
    not g2356(n628 ,n31[0]);
    not g2357(n627 ,n27[1]);
    not g2358(n626 ,n12[4]);
    not g2359(n625 ,n51[6]);
    not g2360(n624 ,n35[0]);
    not g2361(n623 ,n45[3]);
    not g2362(n622 ,n49[5]);
    not g2363(n621 ,n54[7]);
    not g2364(n620 ,n47[0]);
    not g2365(n619 ,n49[7]);
    not g2366(n618 ,n20[2]);
    not g2367(n617 ,n46[4]);
    not g2368(n616 ,n43[2]);
    not g2369(n615 ,n31[4]);
    not g2370(n614 ,n46[7]);
    not g2371(n613 ,n44[2]);
    not g2372(n612 ,n49[2]);
    not g2373(n611 ,n42[2]);
    not g2374(n610 ,n54[3]);
    not g2375(n609 ,n34[3]);
    not g2376(n608 ,n29[5]);
    not g2377(n607 ,n42[7]);
    not g2378(n606 ,n23[4]);
    not g2379(n605 ,n33[4]);
    not g2380(n604 ,n61[3]);
    not g2381(n603 ,n61[7]);
    not g2382(n602 ,n56[4]);
    not g2383(n601 ,n52[0]);
    not g2384(n600 ,n51[0]);
    not g2385(n599 ,n21[0]);
    not g2386(n598 ,n54[6]);
    not g2387(n597 ,n50[0]);
    not g2388(n596 ,n42[3]);
    not g2389(n595 ,n54[5]);
    not g2390(n594 ,n57[1]);
    not g2391(n593 ,n29[7]);
    not g2392(n592 ,n49[0]);
    not g2393(n591 ,n24[3]);
    not g2394(n590 ,n61[6]);
    not g2395(n589 ,n25[5]);
    not g2396(n588 ,n55[5]);
    not g2397(n587 ,n52[3]);
    not g2398(n586 ,n43[5]);
    not g2399(n585 ,n34[6]);
    not g2400(n584 ,n24[0]);
    not g2401(n583 ,n46[0]);
    not g2402(n582 ,n34[0]);
    not g2403(n581 ,n42[1]);
    not g2404(n580 ,n31[7]);
    not g2405(n579 ,n34[5]);
    not g2406(n578 ,n31[2]);
    not g2407(n577 ,n47[6]);
    not g2408(n576 ,n22[3]);
    not g2409(n575 ,n14[1]);
    not g2410(n574 ,n30[7]);
    not g2411(n573 ,n61[2]);
    not g2412(n572 ,n50[2]);
    not g2413(n571 ,n50[3]);
    not g2414(n570 ,n48[0]);
    not g2415(n569 ,n44[1]);
    not g2416(n568 ,n29[6]);
    not g2417(n567 ,n43[3]);
    not g2418(n566 ,n20[3]);
    not g2419(n565 ,n48[1]);
    not g2420(n564 ,n51[2]);
    not g2421(n563 ,n52[6]);
    not g2422(n562 ,n36[0]);
    not g2423(n561 ,n42[6]);
    not g2424(n560 ,n34[2]);
    not g2425(n559 ,n25[0]);
    not g2426(n558 ,n31[6]);
    not g2427(n557 ,n53[5]);
    not g2428(n556 ,n57[7]);
    not g2429(n555 ,n47[3]);
    not g2430(n554 ,n47[1]);
    not g2431(n553 ,n56[6]);
    not g2432(n552 ,n50[1]);
    not g2433(n551 ,n22[5]);
    not g2434(n550 ,n20[1]);
    not g2435(n549 ,n61[4]);
    not g2436(n548 ,n23[2]);
    not g2437(n547 ,n51[3]);
    not g2438(n546 ,n53[6]);
    not g2439(n545 ,n61[1]);
    not g2440(n544 ,n49[1]);
    not g2441(n543 ,n61[0]);
    not g2442(n542 ,n20[11]);
    not g2443(n541 ,n47[2]);
    not g2444(n540 ,n35[2]);
    not g2445(n539 ,n52[1]);
    not g2446(n538 ,n30[1]);
    not g2447(n537 ,n27[5]);
    not g2448(n536 ,n28[6]);
    not g2449(n535 ,n40[5]);
    not g2450(n534 ,n58[0]);
    not g2451(n533 ,n8);
    not g2452(n532 ,n19[2]);
    not g2453(n531 ,n40[1]);
    not g2454(n530 ,n10);
    not g2455(n529 ,n19[1]);
    not g2456(n528 ,n58[2]);
    not g2457(n527 ,n58[3]);
    not g2458(n526 ,n40[3]);
    not g2459(n525 ,n19[3]);
    not g2460(n524 ,n9);
    not g2461(n523 ,n18[1]);
    not g2462(n522 ,n20[0]);
    not g2463(n521 ,n40[8]);
    not g2464(n520 ,n40[4]);
    not g2465(n519 ,n58[1]);
    not g2466(n518 ,n40[9]);
    not g2467(n517 ,n11);
    not g2468(n516 ,n40[10]);
    not g2469(n515 ,n59[3]);
    not g2470(n514 ,n41[1]);
    not g2471(n513 ,n38[0]);
    not g2472(n512 ,n18[0]);
    not g2473(n511 ,n19[4]);
    not g2474(n510 ,n41[0]);
    not g2475(n509 ,n59[2]);
    not g2476(n508 ,n59[1]);
    not g2477(n507 ,n60[1]);
    not g2478(n506 ,n38[2]);
    not g2479(n505 ,n38[3]);
    not g2480(n504 ,n38[1]);
    not g2481(n503 ,n60[2]);
    not g2482(n502 ,n37[0]);
    not g2483(n501 ,n59[0]);
    not g2484(n500 ,n17[0]);
    not g2485(n499 ,n17[1]);
    not g2486(n498 ,n17[2]);
    not g2487(n497 ,n39[0]);
    not g2488(n496 ,n39[2]);
    not g2489(n495 ,n39[7]);
    not g2490(n494 ,n39[5]);
    not g2491(n493 ,n2613);
    not g2492(n492 ,n2637);
    not g2493(n491 ,n2634);
    not g2494(n490 ,n2620);
    not g2495(n489 ,n2628);
    not g2496(n488 ,n2629);
    not g2497(n487 ,n2604);
    not g2498(n486 ,n2636);
    not g2499(n485 ,n2650);
    not g2500(n484 ,n2624);
    not g2501(n483 ,n2649);
    not g2502(n482 ,n2630);
    not g2503(n481 ,n2645);
    not g2504(n480 ,n2633);
    not g2505(n479 ,n2627);
    not g2506(n478 ,n2609);
    not g2507(n477 ,n2598);
    not g2508(n476 ,n2643);
    not g2509(n475 ,n2644);
    not g2510(n474 ,n2648);
    not g2511(n473 ,n2617);
    not g2512(n472 ,n2600);
    not g2513(n471 ,n2610);
    not g2514(n470 ,n2603);
    not g2515(n469 ,n2639);
    not g2516(n468 ,n2640);
    not g2517(n467 ,n2615);
    not g2518(n466 ,n2622);
    not g2519(n465 ,n2608);
    not g2520(n464 ,n2632);
    not g2521(n463 ,n2619);
    not g2522(n462 ,n2616);
    not g2523(n461 ,n2607);
    not g2524(n460 ,n2623);
    not g2525(n459 ,n2635);
    not g2526(n458 ,n2614);
    not g2527(n457 ,n2642);
    not g2528(n456 ,n2625);
    not g2529(n455 ,n2602);
    not g2530(n454 ,n2611);
    not g2531(n453 ,n2605);
    not g2532(n452 ,n2626);
    not g2533(n451 ,n2612);
    not g2534(n450 ,n2599);
    not g2535(n449 ,n2641);
    not g2536(n448 ,n2606);
    not g2537(n447 ,n2651);
    not g2538(n446 ,n2631);
    not g2539(n445 ,n2638);
    not g2540(n444 ,n2601);
    not g2541(n443 ,n50[7]);
    not g2542(n442 ,n24[5]);
    not g2543(n441 ,n30[6]);
    not g2544(n440 ,n23[3]);
    not g2545(n439 ,n34[1]);
    not g2546(n438 ,n22[4]);
    not g2547(n437 ,n54[1]);
    not g2548(n436 ,n48[3]);
    not g2549(n435 ,n55[6]);
    not g2550(n434 ,n36[5]);
    not g2551(n433 ,n36[3]);
    not g2552(n432 ,n21[6]);
    not g2553(n431 ,n20[10]);
    not g2554(n430 ,n47[5]);
    not g2555(n429 ,n52[2]);
    not g2556(n428 ,n30[2]);
    not g2557(n427 ,n35[6]);
    not g2558(n426 ,n25[3]);
    not g2559(n425 ,n52[4]);
    not g2560(n424 ,n61[5]);
    not g2561(n423 ,n20[7]);
    not g2562(n422 ,n21[4]);
    not g2563(n421 ,n57[5]);
    not g2564(n420 ,n12[3]);
    not g2565(n419 ,n50[4]);
    not g2566(n418 ,n21[2]);
    not g2567(n417 ,n46[6]);
    not g2568(n416 ,n57[0]);
    not g2569(n415 ,n32[3]);
    not g2570(n414 ,n51[4]);
    not g2571(n413 ,n26[0]);
    not g2572(n412 ,n26[2]);
    not g2573(n411 ,n45[7]);
    not g2574(n410 ,n32[1]);
    not g2575(n409 ,n32[4]);
    not g2576(n408 ,n28[5]);
    not g2577(n407 ,n57[4]);
    not g2578(n406 ,n33[0]);
    not g2579(n405 ,n53[2]);
    not g2580(n404 ,n45[1]);
    not g2581(n403 ,n26[7]);
    not g2582(n402 ,n43[1]);
    not g2583(n401 ,n57[6]);
    not g2584(n400 ,n27[0]);
    not g2585(n399 ,n36[6]);
    not g2586(n398 ,n24[2]);
    not g2587(n397 ,n48[7]);
    not g2588(n396 ,n35[3]);
    not g2589(n395 ,n56[1]);
    not g2590(n394 ,n49[6]);
    not g2591(n393 ,n28[4]);
    not g2592(n392 ,n44[4]);
    not g2593(n391 ,n48[5]);
    not g2594(n390 ,n12[6]);
    not g2595(n389 ,n21[3]);
    not g2596(n388 ,n48[6]);
    not g2597(n387 ,n56[5]);
    not g2598(n386 ,n22[1]);
    not g2599(n385 ,n28[0]);
    not g2600(n384 ,n22[7]);
    not g2601(n383 ,n31[1]);
    not g2602(n382 ,n25[4]);
    not g2603(n381 ,n53[4]);
    not g2604(n380 ,n30[3]);
    not g2605(n379 ,n36[2]);
    not g2606(n378 ,n27[4]);
    not g2607(n377 ,n42[4]);
    not g2608(n376 ,n12[7]);
    not g2609(n375 ,n36[4]);
    not g2610(n374 ,n44[6]);
    not g2611(n373 ,n51[5]);
    not g2612(n372 ,n26[1]);
    not g2613(n371 ,n44[3]);
    not g2614(n370 ,n55[3]);
    not g2615(n369 ,n42[0]);
    not g2616(n368 ,n46[1]);
    not g2617(n367 ,n22[6]);
    not g2618(n366 ,n56[2]);
    not g2619(n365 ,n55[1]);
    not g2620(n364 ,n22[2]);
    not g2621(n363 ,n48[4]);
    not g2622(n362 ,n33[7]);
    not g2623(n361 ,n26[3]);
    not g2624(n360 ,n42[5]);
    not g2625(n359 ,n20[4]);
    not g2626(n358 ,n28[1]);
    not g2627(n357 ,n36[1]);
    not g2628(n356 ,n55[7]);
    not g2629(n355 ,n56[7]);
    not g2630(n354 ,n24[1]);
    not g2631(n353 ,n56[0]);
    not g2632(n352 ,n30[4]);
    not g2633(n351 ,n31[5]);
    not g2634(n350 ,n23[7]);
    not g2635(n349 ,n24[4]);
    not g2636(n348 ,n21[5]);
    not g2637(n347 ,n55[2]);
    not g2638(n346 ,n32[5]);
    not g2639(n345 ,n49[3]);
    not g2640(n344 ,n23[1]);
    not g2641(n343 ,n48[2]);
    not g2642(n342 ,n50[5]);
    not g2643(n341 ,n52[5]);
    not g2644(n340 ,n50[6]);
    not g2645(n339 ,n34[4]);
    not g2646(n338 ,n45[0]);
    not g2647(n337 ,n23[5]);
    not g2648(n336 ,n45[5]);
    not g2649(n335 ,n33[3]);
    not g2650(n334 ,n35[5]);
    not g2651(n333 ,n45[2]);
    not g2652(n332 ,n29[2]);
    not g2653(n331 ,n30[0]);
    not g2654(n330 ,n12[5]);
    not g2655(n329 ,n32[0]);
    not g2656(n328 ,n2646);
    not g2657(n327 ,n33[6]);
    not g2658(n326 ,n45[4]);
    not g2659(n325 ,n57[3]);
    not g2660(n324 ,n35[4]);
    not g2661(n323 ,n57[2]);
    not g2662(n322 ,n46[5]);
    not g2663(n321 ,n32[6]);
    not g2664(n320 ,n4);
    not g2665(n319 ,n32[2]);
    not g2666(n318 ,n32[7]);
    not g2667(n317 ,n18[2]);
    not g2668(n316 ,n2653);
    not g2669(n315 ,n40[7]);
    not g2670(n314 ,n40[6]);
    not g2671(n313 ,n2654);
    not g2672(n312 ,n40[2]);
    not g2673(n311 ,n40[0]);
    not g2674(n310 ,n41[2]);
    not g2675(n309 ,n37[3]);
    not g2676(n308 ,n62[0]);
    not g2677(n307 ,n62[1]);
    not g2678(n306 ,n60[3]);
    not g2679(n305 ,n2);
    not g2680(n304 ,n58[4]);
    not g2681(n303 ,n37[2]);
    not g2682(n302 ,n37[1]);
    not g2683(n301 ,n60[0]);
    not g2684(n300 ,n2655);
    not g2685(n299 ,n62[2]);
    not g2686(n298 ,n5[7]);
    not g2687(n297 ,n5[2]);
    not g2688(n296 ,n5[6]);
    not g2689(n295 ,n5[0]);
    not g2690(n294 ,n5[4]);
    not g2691(n293 ,n5[3]);
    not g2692(n292 ,n5[5]);
    not g2693(n291 ,n5[1]);
    not g2694(n290 ,n39[4]);
    not g2695(n289 ,n39[3]);
    not g2696(n288 ,n39[6]);
    not g2697(n287 ,n39[1]);
    not g2698(n286 ,n1);
    not g2699(n285 ,n1);
    not g2700(n284 ,n1);
    not g2701(n283 ,n1);
    not g2702(n282 ,n1);
    not g2703(n281 ,n1);
    not g2704(n280 ,n1);
    not g2705(n279 ,n1);
    not g2706(n278 ,n1);
    xor g2707(n2648 ,n19[4] ,n83);
    or g2708(n2649 ,n84 ,n82);
    nor g2709(n84 ,n76 ,n81);
    nor g2710(n83 ,n80 ,n78);
    nor g2711(n82 ,n19[3] ,n79);
    xnor g2712(n2650 ,n19[2] ,n75);
    not g2713(n81 ,n80);
    nor g2714(n80 ,n63 ,n77);
    nor g2715(n79 ,n77 ,n76);
    nor g2716(n78 ,n19[3] ,n76);
    xnor g2717(n2651 ,n19[0] ,n70);
    nor g2718(n77 ,n67 ,n74);
    nor g2719(n76 ,n19[2] ,n72);
    nor g2720(n75 ,n73 ,n71);
    not g2721(n74 ,n73);
    nor g2722(n73 ,n66 ,n69);
    not g2723(n72 ,n71);
    nor g2724(n71 ,n19[0] ,n68);
    xnor g2725(n70 ,n2618 ,n19[1]);
    or g2726(n69 ,n64 ,n2618);
    or g2727(n68 ,n65 ,n19[1]);
    not g2728(n67 ,n19[2]);
    not g2729(n66 ,n19[0]);
    not g2730(n65 ,n2618);
    not g2731(n64 ,n19[1]);
    not g2732(n63 ,n19[3]);
    xor g2733(n2639 ,n58[4] ,n89);
    xor g2734(n2638 ,n58[3] ,n87);
    nor g2735(n89 ,n58[3] ,n88);
    xor g2736(n2637 ,n58[2] ,n85);
    not g2737(n88 ,n87);
    nor g2738(n87 ,n58[2] ,n86);
    xnor g2739(n2636 ,n58[1] ,n58[0]);
    not g2740(n86 ,n85);
    nor g2741(n85 ,n58[1] ,n58[0]);
    or g2742(n2647 ,n91 ,n92);
    or g2743(n92 ,n58[3] ,n90);
    or g2744(n91 ,n58[2] ,n58[0]);
    or g2745(n90 ,n58[4] ,n58[1]);
    or g2746(n2653 ,n94 ,n95);
    or g2747(n95 ,n19[3] ,n93);
    or g2748(n94 ,n19[2] ,n19[0]);
    or g2749(n93 ,n19[4] ,n19[1]);
    or g2750(n2655 ,n40[10] ,n110);
    nor g2751(n110 ,n104 ,n109);
    nor g2752(n109 ,n40[7] ,n108);
    nor g2753(n108 ,n98 ,n107);
    or g2754(n107 ,n100 ,n106);
    nor g2755(n106 ,n102 ,n105);
    or g2756(n105 ,n40[2] ,n103);
    or g2757(n104 ,n101 ,n99);
    nor g2758(n103 ,n96 ,n97);
    or g2759(n102 ,n40[4] ,n40[3]);
    not g2760(n101 ,n40[9]);
    not g2761(n100 ,n40[6]);
    not g2762(n99 ,n40[8]);
    not g2763(n98 ,n40[5]);
    not g2764(n97 ,n40[0]);
    not g2765(n96 ,n40[1]);
    or g2766(n2621 ,n116 ,n125);
    or g2767(n125 ,n20[9] ,n124);
    or g2768(n124 ,n20[12] ,n123);
    nor g2769(n123 ,n118 ,n122);
    nor g2770(n122 ,n20[6] ,n121);
    nor g2771(n121 ,n119 ,n120);
    nor g2772(n120 ,n117 ,n115);
    or g2773(n119 ,n111 ,n113);
    or g2774(n118 ,n112 ,n114);
    or g2775(n117 ,n20[3] ,n20[2]);
    or g2776(n116 ,n20[11] ,n20[10]);
    or g2777(n115 ,n20[1] ,n20[0]);
    not g2778(n114 ,n20[7]);
    not g2779(n113 ,n20[4]);
    not g2780(n112 ,n20[8]);
    not g2781(n111 ,n20[5]);
    or g2782(n2654 ,n132 ,n142);
    or g2783(n142 ,n20[12] ,n141);
    nor g2784(n141 ,n135 ,n140);
    nor g2785(n140 ,n20[7] ,n139);
    nor g2786(n139 ,n131 ,n138);
    or g2787(n138 ,n127 ,n137);
    nor g2788(n137 ,n133 ,n136);
    or g2789(n136 ,n20[2] ,n134);
    or g2790(n135 ,n128 ,n130);
    nor g2791(n134 ,n126 ,n129);
    or g2792(n133 ,n20[4] ,n20[3]);
    or g2793(n132 ,n20[11] ,n20[10]);
    not g2794(n131 ,n20[5]);
    not g2795(n130 ,n20[8]);
    not g2796(n129 ,n20[0]);
    not g2797(n128 ,n20[9]);
    not g2798(n127 ,n20[6]);
    not g2799(n126 ,n20[1]);
    xor g2800(n2600 ,n60[3] ,n150);
    nor g2801(n2599 ,n149 ,n150);
    nor g2802(n150 ,n145 ,n148);
    nor g2803(n149 ,n60[2] ,n147);
    nor g2804(n2598 ,n147 ,n146);
    not g2805(n148 ,n147);
    nor g2806(n147 ,n143 ,n144);
    nor g2807(n146 ,n60[1] ,n60[0]);
    not g2808(n145 ,n60[2]);
    not g2809(n144 ,n60[0]);
    not g2810(n143 ,n60[1]);
    xor g2811(n2643 ,n58[4] ,n162);
    nor g2812(n2642 ,n161 ,n162);
    nor g2813(n162 ,n152 ,n160);
    nor g2814(n161 ,n58[3] ,n159);
    nor g2815(n2641 ,n158 ,n159);
    not g2816(n160 ,n159);
    nor g2817(n159 ,n154 ,n157);
    nor g2818(n158 ,n58[2] ,n156);
    nor g2819(n2640 ,n156 ,n155);
    not g2820(n157 ,n156);
    nor g2821(n156 ,n151 ,n153);
    nor g2822(n155 ,n58[1] ,n58[0]);
    not g2823(n154 ,n58[2]);
    not g2824(n153 ,n58[0]);
    not g2825(n152 ,n58[3]);
    not g2826(n151 ,n58[1]);
    xor g2827(n2603 ,n59[3] ,n170);
    nor g2828(n2602 ,n169 ,n170);
    nor g2829(n170 ,n165 ,n168);
    nor g2830(n169 ,n59[2] ,n167);
    nor g2831(n2601 ,n167 ,n166);
    not g2832(n168 ,n167);
    nor g2833(n167 ,n163 ,n164);
    nor g2834(n166 ,n59[1] ,n59[0]);
    not g2835(n165 ,n59[2]);
    not g2836(n164 ,n59[0]);
    not g2837(n163 ,n59[1]);
    xor g2838(n2635 ,n40[10] ,n206);
    nor g2839(n2634 ,n205 ,n206);
    nor g2840(n206 ,n171 ,n204);
    nor g2841(n205 ,n40[9] ,n203);
    nor g2842(n2633 ,n202 ,n203);
    not g2843(n204 ,n203);
    nor g2844(n203 ,n173 ,n201);
    nor g2845(n202 ,n40[8] ,n200);
    nor g2846(n2632 ,n199 ,n200);
    not g2847(n201 ,n200);
    nor g2848(n200 ,n179 ,n198);
    nor g2849(n199 ,n40[7] ,n197);
    nor g2850(n2631 ,n196 ,n197);
    not g2851(n198 ,n197);
    nor g2852(n197 ,n174 ,n195);
    nor g2853(n196 ,n40[6] ,n194);
    nor g2854(n2630 ,n193 ,n194);
    not g2855(n195 ,n194);
    nor g2856(n194 ,n175 ,n192);
    nor g2857(n193 ,n40[5] ,n191);
    nor g2858(n2629 ,n190 ,n191);
    not g2859(n192 ,n191);
    nor g2860(n191 ,n172 ,n189);
    nor g2861(n190 ,n40[4] ,n188);
    nor g2862(n2628 ,n187 ,n188);
    not g2863(n189 ,n188);
    nor g2864(n188 ,n178 ,n186);
    nor g2865(n187 ,n40[3] ,n185);
    nor g2866(n2627 ,n184 ,n185);
    not g2867(n186 ,n185);
    nor g2868(n185 ,n176 ,n183);
    nor g2869(n184 ,n40[2] ,n182);
    nor g2870(n2626 ,n182 ,n181);
    not g2871(n183 ,n182);
    nor g2872(n182 ,n177 ,n180);
    nor g2873(n181 ,n40[1] ,n40[0]);
    not g2874(n180 ,n40[0]);
    not g2875(n179 ,n40[7]);
    not g2876(n178 ,n40[3]);
    not g2877(n177 ,n40[1]);
    not g2878(n176 ,n40[2]);
    not g2879(n175 ,n40[5]);
    not g2880(n174 ,n40[6]);
    not g2881(n173 ,n40[8]);
    not g2882(n172 ,n40[4]);
    not g2883(n171 ,n40[9]);
    xor g2884(n2645 ,n41[2] ,n210);
    nor g2885(n2644 ,n210 ,n209);
    nor g2886(n210 ,n208 ,n207);
    nor g2887(n209 ,n41[1] ,n41[0]);
    not g2888(n208 ,n41[1]);
    not g2889(n207 ,n41[0]);
    xor g2890(n2606 ,n37[3] ,n218);
    nor g2891(n2605 ,n217 ,n218);
    nor g2892(n218 ,n213 ,n216);
    nor g2893(n217 ,n37[2] ,n215);
    nor g2894(n2604 ,n215 ,n214);
    not g2895(n216 ,n215);
    nor g2896(n215 ,n211 ,n212);
    nor g2897(n214 ,n37[1] ,n37[0]);
    not g2898(n213 ,n37[2]);
    not g2899(n212 ,n37[0]);
    not g2900(n211 ,n37[1]);
    xor g2901(n2617 ,n20[12] ,n262);
    nor g2902(n2616 ,n261 ,n262);
    nor g2903(n262 ,n228 ,n260);
    nor g2904(n261 ,n20[11] ,n259);
    nor g2905(n2615 ,n258 ,n259);
    not g2906(n260 ,n259);
    nor g2907(n259 ,n221 ,n257);
    nor g2908(n258 ,n20[10] ,n256);
    nor g2909(n2614 ,n255 ,n256);
    not g2910(n257 ,n256);
    nor g2911(n256 ,n222 ,n254);
    nor g2912(n255 ,n20[9] ,n253);
    nor g2913(n2625 ,n252 ,n253);
    not g2914(n254 ,n253);
    nor g2915(n253 ,n226 ,n251);
    nor g2916(n252 ,n20[8] ,n250);
    nor g2917(n2613 ,n249 ,n250);
    not g2918(n251 ,n250);
    nor g2919(n250 ,n220 ,n248);
    nor g2920(n249 ,n20[7] ,n247);
    nor g2921(n2624 ,n246 ,n247);
    not g2922(n248 ,n247);
    nor g2923(n247 ,n225 ,n245);
    nor g2924(n246 ,n20[6] ,n244);
    nor g2925(n2612 ,n243 ,n244);
    not g2926(n245 ,n244);
    nor g2927(n244 ,n223 ,n242);
    nor g2928(n243 ,n20[5] ,n241);
    nor g2929(n2623 ,n240 ,n241);
    not g2930(n242 ,n241);
    nor g2931(n241 ,n224 ,n239);
    nor g2932(n240 ,n20[4] ,n238);
    nor g2933(n2611 ,n237 ,n238);
    not g2934(n239 ,n238);
    nor g2935(n238 ,n229 ,n236);
    nor g2936(n237 ,n20[3] ,n235);
    nor g2937(n2622 ,n234 ,n235);
    not g2938(n236 ,n235);
    nor g2939(n235 ,n230 ,n233);
    nor g2940(n234 ,n20[2] ,n232);
    nor g2941(n2610 ,n232 ,n231);
    not g2942(n233 ,n232);
    nor g2943(n232 ,n219 ,n227);
    nor g2944(n231 ,n20[1] ,n20[0]);
    not g2945(n230 ,n20[2]);
    not g2946(n229 ,n20[3]);
    not g2947(n228 ,n20[11]);
    not g2948(n227 ,n20[0]);
    not g2949(n226 ,n20[8]);
    not g2950(n225 ,n20[6]);
    not g2951(n224 ,n20[4]);
    not g2952(n223 ,n20[5]);
    not g2953(n222 ,n20[9]);
    not g2954(n221 ,n20[10]);
    not g2955(n220 ,n20[7]);
    not g2956(n219 ,n20[1]);
    xor g2957(n2620 ,n18[2] ,n266);
    nor g2958(n2619 ,n266 ,n265);
    nor g2959(n266 ,n264 ,n263);
    nor g2960(n265 ,n18[1] ,n18[0]);
    not g2961(n264 ,n18[1]);
    not g2962(n263 ,n18[0]);
    xor g2963(n2609 ,n38[3] ,n274);
    nor g2964(n2608 ,n273 ,n274);
    nor g2965(n274 ,n269 ,n272);
    nor g2966(n273 ,n38[2] ,n271);
    nor g2967(n2607 ,n271 ,n270);
    not g2968(n272 ,n271);
    nor g2969(n271 ,n267 ,n268);
    nor g2970(n270 ,n38[1] ,n38[0]);
    not g2971(n269 ,n38[2]);
    not g2972(n268 ,n38[0]);
    not g2973(n267 ,n38[1]);
    nor g2974(n2652 ,n19[4] ,n277);
    nor g2975(n277 ,n275 ,n276);
    not g2976(n276 ,n19[2]);
    not g2977(n275 ,n19[3]);
    buf g2978(n1326 ,n782);
    not g2979(n881 ,n1);
    buf g2980(n2166 ,n1328);
endmodule
